library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity program_tb is
end entity;

architecture TB of program_tb is
begin
end architecture;
