----------------------------------------------------------------------------
----------------------------------------------------------------------------
--  The Free IP Project
--  VHDL DES Core
--  (c) 1999, The Free IP Project and David Kessner
--
--
--  FREE IP GENERAL PUBLIC LICENSE
--  TERMS AND CONDITIONS FOR USE, COPYING, DISTRIBUTION, AND MODIFICATION
--
--  1.  You may copy and distribute verbatim copies of this core, as long
--      as this file, and the other associated files, remain intact and
--      unmodified.  Modifications are outlined below.  Also, see the
--      import/export warning above for further restrictions on
--      distribution.
--  2.  You may use this core in any way, be it academic, commercial, or
--      military.  Modified or not.
--  3.  Distribution of this core must be free of charge.  Charging is
--      allowed only for value added services.  Value added services
--      would include copying fees, modifications, customizations, and
--      inclusion in other products.
--  4.  If a modified source code is distributed, the original unmodified
--      source code must also be included (or a link to the Free IP web
--      site).  In the modified source code there must be clear
--      identification of the modified version.
--  5.  Visit the Free IP web site for additional information.
--      http://www.free-ip.com
--
----------------------------------------------------------------------------
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library work;

package test_suite is
  component test_rom
    port (addr	:in std_logic_vector (11 downto 0);
          data  :out std_logic_vector (7 downto 0)
         );
  end component;
end test_suite;


------------------------------------------------------------------------------
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library work;
use work.test_suite.all;

entity test_rom is
    port (addr	:in std_logic_vector (11 downto 0);
          data  :out std_logic_vector (7 downto 0)
         );
end test_rom;

architecture arch_test_rom of test_rom is
begin
  process (addr)
  begin
    case addr(11 downto 0) is
      --addrbits 12
      --databits 8
      --varname data
      --little-endian
      --start_of_rom      -- rom2vhdl output.  Tue Jun 20 14:20:58 2000
      when "000000000000" =>  data <= "11101010";  -- 0 = EA
      when "000000000001" =>  data <= "11101010";  -- 1 = EA
      when "000000000010" =>  data <= "11101010";  -- 2 = EA
      when "000000000011" =>  data <= "11101010";  -- 3 = EA
      when "000000000100" =>  data <= "10101001";  -- 4 = A9
      when "000000000101" =>  data <= "00000000";  -- 5 = 0
      when "000000000110" =>  data <= "10000101";  -- 6 = 85
      when "000000000111" =>  data <= "00000100";  -- 7 = 4
      when "000000001000" =>  data <= "10000101";  -- 8 = 85
      when "000000001001" =>  data <= "00000101";  -- 9 = 5
      when "000000001010" =>  data <= "10000101";  -- A = 85
      when "000000001011" =>  data <= "00000110";  -- B = 6
      when "000000001100" =>  data <= "10000101";  -- C = 85
      when "000000001101" =>  data <= "00000111";  -- D = 7
      when "000000001110" =>  data <= "10101001";  -- E = A9
      when "000000001111" =>  data <= "00000000";  -- F = 0
      when "000000010000" =>  data <= "10001101";  -- 10 = 8D
      when "000000010001" =>  data <= "00000001";  -- 11 = 1
      when "000000010010" =>  data <= "10000000";  -- 12 = 80
      when "000000010011" =>  data <= "10101001";  -- 13 = A9
      when "000000010100" =>  data <= "00000001";  -- 14 = 1
      when "000000010101" =>  data <= "10001101";  -- 15 = 8D
      when "000000010110" =>  data <= "00000001";  -- 16 = 1
      when "000000010111" =>  data <= "10000000";  -- 17 = 80
      when "000000011000" =>  data <= "01001100";  -- 18 = 4C
      when "000000011001" =>  data <= "00100000";  -- 19 = 20
      when "000000011010" =>  data <= "11110000";  -- 1A = F0
      when "000000011011" =>  data <= "10101001";  -- 1B = A9
      when "000000011100" =>  data <= "00000000";  -- 1C = 0
      when "000000011101" =>  data <= "01001100";  -- 1D = 4C
      when "000000011110" =>  data <= "01000001";  -- 1E = 41
      when "000000011111" =>  data <= "11111001";  -- 1F = F9
      when "000000100000" =>  data <= "10101001";  -- 20 = A9
      when "000000100001" =>  data <= "00000001";  -- 21 = 1
      when "000000100010" =>  data <= "10001101";  -- 22 = 8D
      when "000000100011" =>  data <= "00000001";  -- 23 = 1
      when "000000100100" =>  data <= "10000000";  -- 24 = 80
      when "000000100101" =>  data <= "10101001";  -- 25 = A9
      when "000000100110" =>  data <= "00000010";  -- 26 = 2
      when "000000100111" =>  data <= "10001101";  -- 27 = 8D
      when "000000101000" =>  data <= "00000001";  -- 28 = 1
      when "000000101001" =>  data <= "10000000";  -- 29 = 80
      when "000000101010" =>  data <= "00011000";  -- 2A = 18
      when "000000101011" =>  data <= "10010000";  -- 2B = 90
      when "000000101100" =>  data <= "00000101";  -- 2C = 5
      when "000000101101" =>  data <= "10101001";  -- 2D = A9
      when "000000101110" =>  data <= "00000001";  -- 2E = 1
      when "000000101111" =>  data <= "01001100";  -- 2F = 4C
      when "000000110000" =>  data <= "01000001";  -- 30 = 41
      when "000000110001" =>  data <= "11111001";  -- 31 = F9
      when "000000110010" =>  data <= "10101001";  -- 32 = A9
      when "000000110011" =>  data <= "00000011";  -- 33 = 3
      when "000000110100" =>  data <= "10001101";  -- 34 = 8D
      when "000000110101" =>  data <= "00000001";  -- 35 = 1
      when "000000110110" =>  data <= "10000000";  -- 36 = 80
      when "000000110111" =>  data <= "00111000";  -- 37 = 38
      when "000000111000" =>  data <= "10010000";  -- 38 = 90
      when "000000111001" =>  data <= "00000011";  -- 39 = 3
      when "000000111010" =>  data <= "01001100";  -- 3A = 4C
      when "000000111011" =>  data <= "01000010";  -- 3B = 42
      when "000000111100" =>  data <= "11110000";  -- 3C = F0
      when "000000111101" =>  data <= "10101001";  -- 3D = A9
      when "000000111110" =>  data <= "00000010";  -- 3E = 2
      when "000000111111" =>  data <= "01001100";  -- 3F = 4C
      when "000001000000" =>  data <= "01000001";  -- 40 = 41
      when "000001000001" =>  data <= "11111001";  -- 41 = F9
      when "000001000010" =>  data <= "10101001";  -- 42 = A9
      when "000001000011" =>  data <= "00000100";  -- 43 = 4
      when "000001000100" =>  data <= "10001101";  -- 44 = 8D
      when "000001000101" =>  data <= "00000001";  -- 45 = 1
      when "000001000110" =>  data <= "10000000";  -- 46 = 80
      when "000001000111" =>  data <= "00111000";  -- 47 = 38
      when "000001001000" =>  data <= "10110000";  -- 48 = B0
      when "000001001001" =>  data <= "00000101";  -- 49 = 5
      when "000001001010" =>  data <= "10101001";  -- 4A = A9
      when "000001001011" =>  data <= "00000001";  -- 4B = 1
      when "000001001100" =>  data <= "01001100";  -- 4C = 4C
      when "000001001101" =>  data <= "01000001";  -- 4D = 41
      when "000001001110" =>  data <= "11111001";  -- 4E = F9
      when "000001001111" =>  data <= "00011000";  -- 4F = 18
      when "000001010000" =>  data <= "10110000";  -- 50 = B0
      when "000001010001" =>  data <= "00000011";  -- 51 = 3
      when "000001010010" =>  data <= "01001100";  -- 52 = 4C
      when "000001010011" =>  data <= "01011010";  -- 53 = 5A
      when "000001010100" =>  data <= "11110000";  -- 54 = F0
      when "000001010101" =>  data <= "10101001";  -- 55 = A9
      when "000001010110" =>  data <= "00000010";  -- 56 = 2
      when "000001010111" =>  data <= "01001100";  -- 57 = 4C
      when "000001011000" =>  data <= "01000001";  -- 58 = 41
      when "000001011001" =>  data <= "11111001";  -- 59 = F9
      when "000001011010" =>  data <= "10101001";  -- 5A = A9
      when "000001011011" =>  data <= "00000101";  -- 5B = 5
      when "000001011100" =>  data <= "10001101";  -- 5C = 8D
      when "000001011101" =>  data <= "00000001";  -- 5D = 1
      when "000001011110" =>  data <= "10000000";  -- 5E = 80
      when "000001011111" =>  data <= "10101001";  -- 5F = A9
      when "000001100000" =>  data <= "00000101";  -- 60 = 5
      when "000001100001" =>  data <= "11001001";  -- 61 = C9
      when "000001100010" =>  data <= "00000100";  -- 62 = 4
      when "000001100011" =>  data <= "11110000";  -- 63 = F0
      when "000001100100" =>  data <= "00000100";  -- 64 = 4
      when "000001100101" =>  data <= "11001001";  -- 65 = C9
      when "000001100110" =>  data <= "00000101";  -- 66 = 5
      when "000001100111" =>  data <= "11110000";  -- 67 = F0
      when "000001101000" =>  data <= "00000101";  -- 68 = 5
      when "000001101001" =>  data <= "10101001";  -- 69 = A9
      when "000001101010" =>  data <= "00000011";  -- 6A = 3
      when "000001101011" =>  data <= "01001100";  -- 6B = 4C
      when "000001101100" =>  data <= "01000001";  -- 6C = 41
      when "000001101101" =>  data <= "11111001";  -- 6D = F9
      when "000001101110" =>  data <= "10101001";  -- 6E = A9
      when "000001101111" =>  data <= "00000110";  -- 6F = 6
      when "000001110000" =>  data <= "10001101";  -- 70 = 8D
      when "000001110001" =>  data <= "00000001";  -- 71 = 1
      when "000001110010" =>  data <= "10000000";  -- 72 = 80
      when "000001110011" =>  data <= "10101001";  -- 73 = A9
      when "000001110100" =>  data <= "11000100";  -- 74 = C4
      when "000001110101" =>  data <= "11001001";  -- 75 = C9
      when "000001110110" =>  data <= "11100100";  -- 76 = E4
      when "000001110111" =>  data <= "11010000";  -- 77 = D0
      when "000001111000" =>  data <= "00000101";  -- 78 = 5
      when "000001111001" =>  data <= "10101001";  -- 79 = A9
      when "000001111010" =>  data <= "00000100";  -- 7A = 4
      when "000001111011" =>  data <= "01001100";  -- 7B = 4C
      when "000001111100" =>  data <= "01000001";  -- 7C = 41
      when "000001111101" =>  data <= "11111001";  -- 7D = F9
      when "000001111110" =>  data <= "11001001";  -- 7E = C9
      when "000001111111" =>  data <= "11000100";  -- 7F = C4
      when "000010000000" =>  data <= "11010000";  -- 80 = D0
      when "000010000001" =>  data <= "00000011";  -- 81 = 3
      when "000010000010" =>  data <= "01001100";  -- 82 = 4C
      when "000010000011" =>  data <= "10001010";  -- 83 = 8A
      when "000010000100" =>  data <= "11110000";  -- 84 = F0
      when "000010000101" =>  data <= "10101001";  -- 85 = A9
      when "000010000110" =>  data <= "00000101";  -- 86 = 5
      when "000010000111" =>  data <= "01001100";  -- 87 = 4C
      when "000010001000" =>  data <= "01000001";  -- 88 = 41
      when "000010001001" =>  data <= "11111001";  -- 89 = F9
      when "000010001010" =>  data <= "10101001";  -- 8A = A9
      when "000010001011" =>  data <= "00000111";  -- 8B = 7
      when "000010001100" =>  data <= "10001101";  -- 8C = 8D
      when "000010001101" =>  data <= "00000001";  -- 8D = 1
      when "000010001110" =>  data <= "10000000";  -- 8E = 80
      when "000010001111" =>  data <= "10100010";  -- 8F = A2
      when "000010010000" =>  data <= "01000010";  -- 90 = 42
      when "000010010001" =>  data <= "11100000";  -- 91 = E0
      when "000010010010" =>  data <= "00110010";  -- 92 = 32
      when "000010010011" =>  data <= "11110000";  -- 93 = F0
      when "000010010100" =>  data <= "00000100";  -- 94 = 4
      when "000010010101" =>  data <= "11100000";  -- 95 = E0
      when "000010010110" =>  data <= "01000010";  -- 96 = 42
      when "000010010111" =>  data <= "11110000";  -- 97 = F0
      when "000010011000" =>  data <= "00000101";  -- 98 = 5
      when "000010011001" =>  data <= "10101001";  -- 99 = A9
      when "000010011010" =>  data <= "00000110";  -- 9A = 6
      when "000010011011" =>  data <= "01001100";  -- 9B = 4C
      when "000010011100" =>  data <= "01000001";  -- 9C = 41
      when "000010011101" =>  data <= "11111001";  -- 9D = F9
      when "000010011110" =>  data <= "10101001";  -- 9E = A9
      when "000010011111" =>  data <= "00001000";  -- 9F = 8
      when "000010100000" =>  data <= "10001101";  -- A0 = 8D
      when "000010100001" =>  data <= "00000001";  -- A1 = 1
      when "000010100010" =>  data <= "10000000";  -- A2 = 80
      when "000010100011" =>  data <= "10100000";  -- A3 = A0
      when "000010100100" =>  data <= "11000011";  -- A4 = C3
      when "000010100101" =>  data <= "11000000";  -- A5 = C0
      when "000010100110" =>  data <= "11010011";  -- A6 = D3
      when "000010100111" =>  data <= "11110000";  -- A7 = F0
      when "000010101000" =>  data <= "00000100";  -- A8 = 4
      when "000010101001" =>  data <= "11000000";  -- A9 = C0
      when "000010101010" =>  data <= "11000011";  -- AA = C3
      when "000010101011" =>  data <= "11110000";  -- AB = F0
      when "000010101100" =>  data <= "00000101";  -- AC = 5
      when "000010101101" =>  data <= "10101001";  -- AD = A9
      when "000010101110" =>  data <= "00000111";  -- AE = 7
      when "000010101111" =>  data <= "01001100";  -- AF = 4C
      when "000010110000" =>  data <= "01000001";  -- B0 = 41
      when "000010110001" =>  data <= "11111001";  -- B1 = F9
      when "000010110010" =>  data <= "10101001";  -- B2 = A9
      when "000010110011" =>  data <= "00001001";  -- B3 = 9
      when "000010110100" =>  data <= "10001101";  -- B4 = 8D
      when "000010110101" =>  data <= "00000001";  -- B5 = 1
      when "000010110110" =>  data <= "10000000";  -- B6 = 80
      when "000010110111" =>  data <= "10100010";  -- B7 = A2
      when "000010111000" =>  data <= "00000000";  -- B8 = 0
      when "000010111001" =>  data <= "11001010";  -- B9 = CA
      when "000010111010" =>  data <= "11100000";  -- BA = E0
      when "000010111011" =>  data <= "11111111";  -- BB = FF
      when "000010111100" =>  data <= "11110000";  -- BC = F0
      when "000010111101" =>  data <= "00000101";  -- BD = 5
      when "000010111110" =>  data <= "10101001";  -- BE = A9
      when "000010111111" =>  data <= "00001000";  -- BF = 8
      when "000011000000" =>  data <= "01001100";  -- C0 = 4C
      when "000011000001" =>  data <= "01000001";  -- C1 = 41
      when "000011000010" =>  data <= "11111001";  -- C2 = F9
      when "000011000011" =>  data <= "10101001";  -- C3 = A9
      when "000011000100" =>  data <= "00001010";  -- C4 = A
      when "000011000101" =>  data <= "10001101";  -- C5 = 8D
      when "000011000110" =>  data <= "00000001";  -- C6 = 1
      when "000011000111" =>  data <= "10000000";  -- C7 = 80
      when "000011001000" =>  data <= "10100000";  -- C8 = A0
      when "000011001001" =>  data <= "00000000";  -- C9 = 0
      when "000011001010" =>  data <= "10001000";  -- CA = 88
      when "000011001011" =>  data <= "11000000";  -- CB = C0
      when "000011001100" =>  data <= "11111111";  -- CC = FF
      when "000011001101" =>  data <= "11110000";  -- CD = F0
      when "000011001110" =>  data <= "00000101";  -- CE = 5
      when "000011001111" =>  data <= "10101001";  -- CF = A9
      when "000011010000" =>  data <= "00001001";  -- D0 = 9
      when "000011010001" =>  data <= "01001100";  -- D1 = 4C
      when "000011010010" =>  data <= "01000001";  -- D2 = 41
      when "000011010011" =>  data <= "11111001";  -- D3 = F9
      when "000011010100" =>  data <= "10101001";  -- D4 = A9
      when "000011010101" =>  data <= "00001011";  -- D5 = B
      when "000011010110" =>  data <= "10001101";  -- D6 = 8D
      when "000011010111" =>  data <= "00000001";  -- D7 = 1
      when "000011011000" =>  data <= "10000000";  -- D8 = 80
      when "000011011001" =>  data <= "10100010";  -- D9 = A2
      when "000011011010" =>  data <= "00001111";  -- DA = F
      when "000011011011" =>  data <= "11101000";  -- DB = E8
      when "000011011100" =>  data <= "11100000";  -- DC = E0
      when "000011011101" =>  data <= "00010000";  -- DD = 10
      when "000011011110" =>  data <= "11110000";  -- DE = F0
      when "000011011111" =>  data <= "00000101";  -- DF = 5
      when "000011100000" =>  data <= "10101001";  -- E0 = A9
      when "000011100001" =>  data <= "00010000";  -- E1 = 10
      when "000011100010" =>  data <= "01001100";  -- E2 = 4C
      when "000011100011" =>  data <= "01000001";  -- E3 = 41
      when "000011100100" =>  data <= "11111001";  -- E4 = F9
      when "000011100101" =>  data <= "10101001";  -- E5 = A9
      when "000011100110" =>  data <= "00001100";  -- E6 = C
      when "000011100111" =>  data <= "10001101";  -- E7 = 8D
      when "000011101000" =>  data <= "00000001";  -- E8 = 1
      when "000011101001" =>  data <= "10000000";  -- E9 = 80
      when "000011101010" =>  data <= "10100000";  -- EA = A0
      when "000011101011" =>  data <= "01111111";  -- EB = 7F
      when "000011101100" =>  data <= "11001000";  -- EC = C8
      when "000011101101" =>  data <= "11000000";  -- ED = C0
      when "000011101110" =>  data <= "10000000";  -- EE = 80
      when "000011101111" =>  data <= "11110000";  -- EF = F0
      when "000011110000" =>  data <= "00000101";  -- F0 = 5
      when "000011110001" =>  data <= "10101001";  -- F1 = A9
      when "000011110010" =>  data <= "00010001";  -- F2 = 11
      when "000011110011" =>  data <= "01001100";  -- F3 = 4C
      when "000011110100" =>  data <= "01000001";  -- F4 = 41
      when "000011110101" =>  data <= "11111001";  -- F5 = F9
      when "000011110110" =>  data <= "10101001";  -- F6 = A9
      when "000011110111" =>  data <= "00001101";  -- F7 = D
      when "000011111000" =>  data <= "10001101";  -- F8 = 8D
      when "000011111001" =>  data <= "00000001";  -- F9 = 1
      when "000011111010" =>  data <= "10000000";  -- FA = 80
      when "000011111011" =>  data <= "10101001";  -- FB = A9
      when "000011111100" =>  data <= "11101101";  -- FC = ED
      when "000011111101" =>  data <= "00100000";  -- FD = 20
      when "000011111110" =>  data <= "00001001";  -- FE = 9
      when "000011111111" =>  data <= "11110001";  -- FF = F1
      when "000100000000" =>  data <= "11001001";  -- 100 = C9
      when "000100000001" =>  data <= "01000010";  -- 101 = 42
      when "000100000010" =>  data <= "11110000";  -- 102 = F0
      when "000100000011" =>  data <= "00001000";  -- 103 = 8
      when "000100000100" =>  data <= "10101001";  -- 104 = A9
      when "000100000101" =>  data <= "00010010";  -- 105 = 12
      when "000100000110" =>  data <= "01001100";  -- 106 = 4C
      when "000100000111" =>  data <= "01000001";  -- 107 = 41
      when "000100001000" =>  data <= "11111001";  -- 108 = F9
      when "000100001001" =>  data <= "10101001";  -- 109 = A9
      when "000100001010" =>  data <= "01000010";  -- 10A = 42
      when "000100001011" =>  data <= "01100000";  -- 10B = 60
      when "000100001100" =>  data <= "10101001";  -- 10C = A9
      when "000100001101" =>  data <= "00001110";  -- 10D = E
      when "000100001110" =>  data <= "10001101";  -- 10E = 8D
      when "000100001111" =>  data <= "00000001";  -- 10F = 1
      when "000100010000" =>  data <= "10000000";  -- 110 = 80
      when "000100010001" =>  data <= "10101001";  -- 111 = A9
      when "000100010010" =>  data <= "00110101";  -- 112 = 35
      when "000100010011" =>  data <= "10101010";  -- 113 = AA
      when "000100010100" =>  data <= "11100000";  -- 114 = E0
      when "000100010101" =>  data <= "00110101";  -- 115 = 35
      when "000100010110" =>  data <= "11110000";  -- 116 = F0
      when "000100010111" =>  data <= "00000101";  -- 117 = 5
      when "000100011000" =>  data <= "10101001";  -- 118 = A9
      when "000100011001" =>  data <= "00010010";  -- 119 = 12
      when "000100011010" =>  data <= "01001100";  -- 11A = 4C
      when "000100011011" =>  data <= "01000001";  -- 11B = 41
      when "000100011100" =>  data <= "11111001";  -- 11C = F9
      when "000100011101" =>  data <= "10101001";  -- 11D = A9
      when "000100011110" =>  data <= "00001111";  -- 11E = F
      when "000100011111" =>  data <= "10001101";  -- 11F = 8D
      when "000100100000" =>  data <= "00000001";  -- 120 = 1
      when "000100100001" =>  data <= "10000000";  -- 121 = 80
      when "000100100010" =>  data <= "10101001";  -- 122 = A9
      when "000100100011" =>  data <= "01110110";  -- 123 = 76
      when "000100100100" =>  data <= "10101000";  -- 124 = A8
      when "000100100101" =>  data <= "11000000";  -- 125 = C0
      when "000100100110" =>  data <= "01110110";  -- 126 = 76
      when "000100100111" =>  data <= "11110000";  -- 127 = F0
      when "000100101000" =>  data <= "00000101";  -- 128 = 5
      when "000100101001" =>  data <= "10101001";  -- 129 = A9
      when "000100101010" =>  data <= "00010011";  -- 12A = 13
      when "000100101011" =>  data <= "01001100";  -- 12B = 4C
      when "000100101100" =>  data <= "01000001";  -- 12C = 41
      when "000100101101" =>  data <= "11111001";  -- 12D = F9
      when "000100101110" =>  data <= "10101001";  -- 12E = A9
      when "000100101111" =>  data <= "00010000";  -- 12F = 10
      when "000100110000" =>  data <= "10001101";  -- 130 = 8D
      when "000100110001" =>  data <= "00000001";  -- 131 = 1
      when "000100110010" =>  data <= "10000000";  -- 132 = 80
      when "000100110011" =>  data <= "10100010";  -- 133 = A2
      when "000100110100" =>  data <= "01010010";  -- 134 = 52
      when "000100110101" =>  data <= "10001010";  -- 135 = 8A
      when "000100110110" =>  data <= "11001001";  -- 136 = C9
      when "000100110111" =>  data <= "01010010";  -- 137 = 52
      when "000100111000" =>  data <= "11110000";  -- 138 = F0
      when "000100111001" =>  data <= "00000101";  -- 139 = 5
      when "000100111010" =>  data <= "10101001";  -- 13A = A9
      when "000100111011" =>  data <= "00010100";  -- 13B = 14
      when "000100111100" =>  data <= "01001100";  -- 13C = 4C
      when "000100111101" =>  data <= "01000001";  -- 13D = 41
      when "000100111110" =>  data <= "11111001";  -- 13E = F9
      when "000100111111" =>  data <= "10101001";  -- 13F = A9
      when "000101000000" =>  data <= "00010001";  -- 140 = 11
      when "000101000001" =>  data <= "10001101";  -- 141 = 8D
      when "000101000010" =>  data <= "00000001";  -- 142 = 1
      when "000101000011" =>  data <= "10000000";  -- 143 = 80
      when "000101000100" =>  data <= "10100000";  -- 144 = A0
      when "000101000101" =>  data <= "01010010";  -- 145 = 52
      when "000101000110" =>  data <= "10011000";  -- 146 = 98
      when "000101000111" =>  data <= "11001001";  -- 147 = C9
      when "000101001000" =>  data <= "01010010";  -- 148 = 52
      when "000101001001" =>  data <= "11110000";  -- 149 = F0
      when "000101001010" =>  data <= "00000101";  -- 14A = 5
      when "000101001011" =>  data <= "10101001";  -- 14B = A9
      when "000101001100" =>  data <= "00010101";  -- 14C = 15
      when "000101001101" =>  data <= "01001100";  -- 14D = 4C
      when "000101001110" =>  data <= "01000001";  -- 14E = 41
      when "000101001111" =>  data <= "11111001";  -- 14F = F9
      when "000101010000" =>  data <= "10101001";  -- 150 = A9
      when "000101010001" =>  data <= "00010010";  -- 151 = 12
      when "000101010010" =>  data <= "10001101";  -- 152 = 8D
      when "000101010011" =>  data <= "00000001";  -- 153 = 1
      when "000101010100" =>  data <= "10000000";  -- 154 = 80
      when "000101010101" =>  data <= "00011000";  -- 155 = 18
      when "000101010110" =>  data <= "10101001";  -- 156 = A9
      when "000101010111" =>  data <= "00100011";  -- 157 = 23
      when "000101011000" =>  data <= "01101001";  -- 158 = 69
      when "000101011001" =>  data <= "01000101";  -- 159 = 45
      when "000101011010" =>  data <= "11001001";  -- 15A = C9
      when "000101011011" =>  data <= "01101000";  -- 15B = 68
      when "000101011100" =>  data <= "11110000";  -- 15C = F0
      when "000101011101" =>  data <= "00000101";  -- 15D = 5
      when "000101011110" =>  data <= "10101001";  -- 15E = A9
      when "000101011111" =>  data <= "00010110";  -- 15F = 16
      when "000101100000" =>  data <= "01001100";  -- 160 = 4C
      when "000101100001" =>  data <= "01000001";  -- 161 = 41
      when "000101100010" =>  data <= "11111001";  -- 162 = F9
      when "000101100011" =>  data <= "00111000";  -- 163 = 38
      when "000101100100" =>  data <= "10101001";  -- 164 = A9
      when "000101100101" =>  data <= "01000010";  -- 165 = 42
      when "000101100110" =>  data <= "01101001";  -- 166 = 69
      when "000101100111" =>  data <= "01100011";  -- 167 = 63
      when "000101101000" =>  data <= "11001001";  -- 168 = C9
      when "000101101001" =>  data <= "10100110";  -- 169 = A6
      when "000101101010" =>  data <= "11110000";  -- 16A = F0
      when "000101101011" =>  data <= "00000101";  -- 16B = 5
      when "000101101100" =>  data <= "10101001";  -- 16C = A9
      when "000101101101" =>  data <= "00010111";  -- 16D = 17
      when "000101101110" =>  data <= "01001100";  -- 16E = 4C
      when "000101101111" =>  data <= "01000001";  -- 16F = 41
      when "000101110000" =>  data <= "11111001";  -- 170 = F9
      when "000101110001" =>  data <= "10101001";  -- 171 = A9
      when "000101110010" =>  data <= "00010011";  -- 172 = 13
      when "000101110011" =>  data <= "10001101";  -- 173 = 8D
      when "000101110100" =>  data <= "00000001";  -- 174 = 1
      when "000101110101" =>  data <= "10000000";  -- 175 = 80
      when "000101110110" =>  data <= "10101001";  -- 176 = A9
      when "000101110111" =>  data <= "00110110";  -- 177 = 36
      when "000101111000" =>  data <= "00101001";  -- 178 = 29
      when "000101111001" =>  data <= "11110000";  -- 179 = F0
      when "000101111010" =>  data <= "11001001";  -- 17A = C9
      when "000101111011" =>  data <= "00110000";  -- 17B = 30
      when "000101111100" =>  data <= "11110000";  -- 17C = F0
      when "000101111101" =>  data <= "00000101";  -- 17D = 5
      when "000101111110" =>  data <= "10101001";  -- 17E = A9
      when "000101111111" =>  data <= "00011000";  -- 17F = 18
      when "000110000000" =>  data <= "01001100";  -- 180 = 4C
      when "000110000001" =>  data <= "01000001";  -- 181 = 41
      when "000110000010" =>  data <= "11111001";  -- 182 = F9
      when "000110000011" =>  data <= "10101001";  -- 183 = A9
      when "000110000100" =>  data <= "00010100";  -- 184 = 14
      when "000110000101" =>  data <= "10001101";  -- 185 = 8D
      when "000110000110" =>  data <= "00000001";  -- 186 = 1
      when "000110000111" =>  data <= "10000000";  -- 187 = 80
      when "000110001000" =>  data <= "00011000";  -- 188 = 18
      when "000110001001" =>  data <= "10101001";  -- 189 = A9
      when "000110001010" =>  data <= "00110110";  -- 18A = 36
      when "000110001011" =>  data <= "00001010";  -- 18B = A
      when "000110001100" =>  data <= "11001001";  -- 18C = C9
      when "000110001101" =>  data <= "01101100";  -- 18D = 6C
      when "000110001110" =>  data <= "11110000";  -- 18E = F0
      when "000110001111" =>  data <= "00000101";  -- 18F = 5
      when "000110010000" =>  data <= "10101001";  -- 190 = A9
      when "000110010001" =>  data <= "00011001";  -- 191 = 19
      when "000110010010" =>  data <= "01001100";  -- 192 = 4C
      when "000110010011" =>  data <= "01000001";  -- 193 = 41
      when "000110010100" =>  data <= "11111001";  -- 194 = F9
      when "000110010101" =>  data <= "10101001";  -- 195 = A9
      when "000110010110" =>  data <= "00010101";  -- 196 = 15
      when "000110010111" =>  data <= "10001101";  -- 197 = 8D
      when "000110011000" =>  data <= "00000001";  -- 198 = 1
      when "000110011001" =>  data <= "10000000";  -- 199 = 80
      when "000110011010" =>  data <= "10101001";  -- 19A = A9
      when "000110011011" =>  data <= "10001001";  -- 19B = 89
      when "000110011100" =>  data <= "01001001";  -- 19C = 49
      when "000110011101" =>  data <= "10010110";  -- 19D = 96
      when "000110011110" =>  data <= "11001001";  -- 19E = C9
      when "000110011111" =>  data <= "00011111";  -- 19F = 1F
      when "000110100000" =>  data <= "11110000";  -- 1A0 = F0
      when "000110100001" =>  data <= "00000101";  -- 1A1 = 5
      when "000110100010" =>  data <= "10101001";  -- 1A2 = A9
      when "000110100011" =>  data <= "00100000";  -- 1A3 = 20
      when "000110100100" =>  data <= "01001100";  -- 1A4 = 4C
      when "000110100101" =>  data <= "01000001";  -- 1A5 = 41
      when "000110100110" =>  data <= "11111001";  -- 1A6 = F9
      when "000110100111" =>  data <= "10101001";  -- 1A7 = A9
      when "000110101000" =>  data <= "00010110";  -- 1A8 = 16
      when "000110101001" =>  data <= "10001101";  -- 1A9 = 8D
      when "000110101010" =>  data <= "00000001";  -- 1AA = 1
      when "000110101011" =>  data <= "10000000";  -- 1AB = 80
      when "000110101100" =>  data <= "00011000";  -- 1AC = 18
      when "000110101101" =>  data <= "10101001";  -- 1AD = A9
      when "000110101110" =>  data <= "01010010";  -- 1AE = 52
      when "000110101111" =>  data <= "01001010";  -- 1AF = 4A
      when "000110110000" =>  data <= "11001001";  -- 1B0 = C9
      when "000110110001" =>  data <= "00101001";  -- 1B1 = 29
      when "000110110010" =>  data <= "11110000";  -- 1B2 = F0
      when "000110110011" =>  data <= "00000101";  -- 1B3 = 5
      when "000110110100" =>  data <= "10101001";  -- 1B4 = A9
      when "000110110101" =>  data <= "00100001";  -- 1B5 = 21
      when "000110110110" =>  data <= "01001100";  -- 1B6 = 4C
      when "000110110111" =>  data <= "01000001";  -- 1B7 = 41
      when "000110111000" =>  data <= "11111001";  -- 1B8 = F9
      when "000110111001" =>  data <= "10101001";  -- 1B9 = A9
      when "000110111010" =>  data <= "00010111";  -- 1BA = 17
      when "000110111011" =>  data <= "10001101";  -- 1BB = 8D
      when "000110111100" =>  data <= "00000001";  -- 1BC = 1
      when "000110111101" =>  data <= "10000000";  -- 1BD = 80
      when "000110111110" =>  data <= "10101001";  -- 1BE = A9
      when "000110111111" =>  data <= "10110110";  -- 1BF = B6
      when "000111000000" =>  data <= "00001001";  -- 1C0 = 9
      when "000111000001" =>  data <= "01001101";  -- 1C1 = 4D
      when "000111000010" =>  data <= "11001001";  -- 1C2 = C9
      when "000111000011" =>  data <= "11111111";  -- 1C3 = FF
      when "000111000100" =>  data <= "11110000";  -- 1C4 = F0
      when "000111000101" =>  data <= "00000101";  -- 1C5 = 5
      when "000111000110" =>  data <= "10101001";  -- 1C6 = A9
      when "000111000111" =>  data <= "00100010";  -- 1C7 = 22
      when "000111001000" =>  data <= "01001100";  -- 1C8 = 4C
      when "000111001001" =>  data <= "01000001";  -- 1C9 = 41
      when "000111001010" =>  data <= "11111001";  -- 1CA = F9
      when "000111001011" =>  data <= "10101001";  -- 1CB = A9
      when "000111001100" =>  data <= "00011000";  -- 1CC = 18
      when "000111001101" =>  data <= "10001101";  -- 1CD = 8D
      when "000111001110" =>  data <= "00000001";  -- 1CE = 1
      when "000111001111" =>  data <= "10000000";  -- 1CF = 80
      when "000111010000" =>  data <= "00011000";  -- 1D0 = 18
      when "000111010001" =>  data <= "10101001";  -- 1D1 = A9
      when "000111010010" =>  data <= "00100011";  -- 1D2 = 23
      when "000111010011" =>  data <= "00101010";  -- 1D3 = 2A
      when "000111010100" =>  data <= "11001001";  -- 1D4 = C9
      when "000111010101" =>  data <= "01000110";  -- 1D5 = 46
      when "000111010110" =>  data <= "11110000";  -- 1D6 = F0
      when "000111010111" =>  data <= "00000101";  -- 1D7 = 5
      when "000111011000" =>  data <= "10101001";  -- 1D8 = A9
      when "000111011001" =>  data <= "00100011";  -- 1D9 = 23
      when "000111011010" =>  data <= "01001100";  -- 1DA = 4C
      when "000111011011" =>  data <= "01000001";  -- 1DB = 41
      when "000111011100" =>  data <= "11111001";  -- 1DC = F9
      when "000111011101" =>  data <= "00111000";  -- 1DD = 38
      when "000111011110" =>  data <= "10101001";  -- 1DE = A9
      when "000111011111" =>  data <= "01000010";  -- 1DF = 42
      when "000111100000" =>  data <= "00101010";  -- 1E0 = 2A
      when "000111100001" =>  data <= "11001001";  -- 1E1 = C9
      when "000111100010" =>  data <= "10000101";  -- 1E2 = 85
      when "000111100011" =>  data <= "11110000";  -- 1E3 = F0
      when "000111100100" =>  data <= "00000101";  -- 1E4 = 5
      when "000111100101" =>  data <= "10101001";  -- 1E5 = A9
      when "000111100110" =>  data <= "00100100";  -- 1E6 = 24
      when "000111100111" =>  data <= "01001100";  -- 1E7 = 4C
      when "000111101000" =>  data <= "01000001";  -- 1E8 = 41
      when "000111101001" =>  data <= "11111001";  -- 1E9 = F9
      when "000111101010" =>  data <= "10101001";  -- 1EA = A9
      when "000111101011" =>  data <= "00011001";  -- 1EB = 19
      when "000111101100" =>  data <= "10001101";  -- 1EC = 8D
      when "000111101101" =>  data <= "00000001";  -- 1ED = 1
      when "000111101110" =>  data <= "10000000";  -- 1EE = 80
      when "000111101111" =>  data <= "00011000";  -- 1EF = 18
      when "000111110000" =>  data <= "10101001";  -- 1F0 = A9
      when "000111110001" =>  data <= "00100011";  -- 1F1 = 23
      when "000111110010" =>  data <= "01101010";  -- 1F2 = 6A
      when "000111110011" =>  data <= "11001001";  -- 1F3 = C9
      when "000111110100" =>  data <= "00010001";  -- 1F4 = 11
      when "000111110101" =>  data <= "11110000";  -- 1F5 = F0
      when "000111110110" =>  data <= "00000101";  -- 1F6 = 5
      when "000111110111" =>  data <= "10101001";  -- 1F7 = A9
      when "000111111000" =>  data <= "00100101";  -- 1F8 = 25
      when "000111111001" =>  data <= "01001100";  -- 1F9 = 4C
      when "000111111010" =>  data <= "01000001";  -- 1FA = 41
      when "000111111011" =>  data <= "11111001";  -- 1FB = F9
      when "000111111100" =>  data <= "00111000";  -- 1FC = 38
      when "000111111101" =>  data <= "10101001";  -- 1FD = A9
      when "000111111110" =>  data <= "01000010";  -- 1FE = 42
      when "000111111111" =>  data <= "01101010";  -- 1FF = 6A
      when "001000000000" =>  data <= "11001001";  -- 200 = C9
      when "001000000001" =>  data <= "10100001";  -- 201 = A1
      when "001000000010" =>  data <= "11110000";  -- 202 = F0
      when "001000000011" =>  data <= "00000101";  -- 203 = 5
      when "001000000100" =>  data <= "10101001";  -- 204 = A9
      when "001000000101" =>  data <= "00100110";  -- 205 = 26
      when "001000000110" =>  data <= "01001100";  -- 206 = 4C
      when "001000000111" =>  data <= "01000001";  -- 207 = 41
      when "001000001000" =>  data <= "11111001";  -- 208 = F9
      when "001000001001" =>  data <= "10101001";  -- 209 = A9
      when "001000001010" =>  data <= "00100000";  -- 20A = 20
      when "001000001011" =>  data <= "10001101";  -- 20B = 8D
      when "001000001100" =>  data <= "00000001";  -- 20C = 1
      when "001000001101" =>  data <= "10000000";  -- 20D = 80
      when "001000001110" =>  data <= "00111000";  -- 20E = 38
      when "001000001111" =>  data <= "10101001";  -- 20F = A9
      when "001000010000" =>  data <= "10000110";  -- 210 = 86
      when "001000010001" =>  data <= "11101001";  -- 211 = E9
      when "001000010010" =>  data <= "01000101";  -- 212 = 45
      when "001000010011" =>  data <= "11001001";  -- 213 = C9
      when "001000010100" =>  data <= "01000001";  -- 214 = 41
      when "001000010101" =>  data <= "11110000";  -- 215 = F0
      when "001000010110" =>  data <= "00000101";  -- 216 = 5
      when "001000010111" =>  data <= "10101001";  -- 217 = A9
      when "001000011000" =>  data <= "00100111";  -- 218 = 27
      when "001000011001" =>  data <= "01001100";  -- 219 = 4C
      when "001000011010" =>  data <= "01000001";  -- 21A = 41
      when "001000011011" =>  data <= "11111001";  -- 21B = F9
      when "001000011100" =>  data <= "00011000";  -- 21C = 18
      when "001000011101" =>  data <= "10101001";  -- 21D = A9
      when "001000011110" =>  data <= "10001001";  -- 21E = 89
      when "001000011111" =>  data <= "11101001";  -- 21F = E9
      when "001000100000" =>  data <= "00100011";  -- 220 = 23
      when "001000100001" =>  data <= "11001001";  -- 221 = C9
      when "001000100010" =>  data <= "01100101";  -- 222 = 65
      when "001000100011" =>  data <= "11110000";  -- 223 = F0
      when "001000100100" =>  data <= "00000101";  -- 224 = 5
      when "001000100101" =>  data <= "10101001";  -- 225 = A9
      when "001000100110" =>  data <= "00101000";  -- 226 = 28
      when "001000100111" =>  data <= "01001100";  -- 227 = 4C
      when "001000101000" =>  data <= "01000001";  -- 228 = 41
      when "001000101001" =>  data <= "11111001";  -- 229 = F9
      when "001000101010" =>  data <= "10101001";  -- 22A = A9
      when "001000101011" =>  data <= "00100001";  -- 22B = 21
      when "001000101100" =>  data <= "10001101";  -- 22C = 8D
      when "001000101101" =>  data <= "00000001";  -- 22D = 1
      when "001000101110" =>  data <= "10000000";  -- 22E = 80
      when "001000101111" =>  data <= "10101001";  -- 22F = A9
      when "001000110000" =>  data <= "01000010";  -- 230 = 42
      when "001000110001" =>  data <= "10001101";  -- 231 = 8D
      when "001000110010" =>  data <= "00000000";  -- 232 = 0
      when "001000110011" =>  data <= "00000010";  -- 233 = 2
      when "001000110100" =>  data <= "10101001";  -- 234 = A9
      when "001000110101" =>  data <= "10011111";  -- 235 = 9F
      when "001000110110" =>  data <= "10001101";  -- 236 = 8D
      when "001000110111" =>  data <= "00000001";  -- 237 = 1
      when "001000111000" =>  data <= "00000010";  -- 238 = 2
      when "001000111001" =>  data <= "10101101";  -- 239 = AD
      when "001000111010" =>  data <= "00000000";  -- 23A = 0
      when "001000111011" =>  data <= "00000010";  -- 23B = 2
      when "001000111100" =>  data <= "11001001";  -- 23C = C9
      when "001000111101" =>  data <= "01000010";  -- 23D = 42
      when "001000111110" =>  data <= "11110000";  -- 23E = F0
      when "001000111111" =>  data <= "00000101";  -- 23F = 5
      when "001001000000" =>  data <= "10101001";  -- 240 = A9
      when "001001000001" =>  data <= "00101001";  -- 241 = 29
      when "001001000010" =>  data <= "01001100";  -- 242 = 4C
      when "001001000011" =>  data <= "01000001";  -- 243 = 41
      when "001001000100" =>  data <= "11111001";  -- 244 = F9
      when "001001000101" =>  data <= "10101101";  -- 245 = AD
      when "001001000110" =>  data <= "00000001";  -- 246 = 1
      when "001001000111" =>  data <= "00000010";  -- 247 = 2
      when "001001001000" =>  data <= "11001001";  -- 248 = C9
      when "001001001001" =>  data <= "10011111";  -- 249 = 9F
      when "001001001010" =>  data <= "11110000";  -- 24A = F0
      when "001001001011" =>  data <= "00000101";  -- 24B = 5
      when "001001001100" =>  data <= "10101001";  -- 24C = A9
      when "001001001101" =>  data <= "00110000";  -- 24D = 30
      when "001001001110" =>  data <= "01001100";  -- 24E = 4C
      when "001001001111" =>  data <= "01000001";  -- 24F = 41
      when "001001010000" =>  data <= "11111001";  -- 250 = F9
      when "001001010001" =>  data <= "10101001";  -- 251 = A9
      when "001001010010" =>  data <= "00100010";  -- 252 = 22
      when "001001010011" =>  data <= "10001101";  -- 253 = 8D
      when "001001010100" =>  data <= "00000001";  -- 254 = 1
      when "001001010101" =>  data <= "10000000";  -- 255 = 80
      when "001001010110" =>  data <= "10101001";  -- 256 = A9
      when "001001010111" =>  data <= "10010100";  -- 257 = 94
      when "001001011000" =>  data <= "10001101";  -- 258 = 8D
      when "001001011001" =>  data <= "00000001";  -- 259 = 1
      when "001001011010" =>  data <= "00000010";  -- 25A = 2
      when "001001011011" =>  data <= "10101001";  -- 25B = A9
      when "001001011100" =>  data <= "01000001";  -- 25C = 41
      when "001001011101" =>  data <= "10001101";  -- 25D = 8D
      when "001001011110" =>  data <= "00000000";  -- 25E = 0
      when "001001011111" =>  data <= "00000010";  -- 25F = 2
      when "001001100000" =>  data <= "10101001";  -- 260 = A9
      when "001001100001" =>  data <= "01010011";  -- 261 = 53
      when "001001100010" =>  data <= "00011000";  -- 262 = 18
      when "001001100011" =>  data <= "01101101";  -- 263 = 6D
      when "001001100100" =>  data <= "00000000";  -- 264 = 0
      when "001001100101" =>  data <= "00000010";  -- 265 = 2
      when "001001100110" =>  data <= "11001101";  -- 266 = CD
      when "001001100111" =>  data <= "00000001";  -- 267 = 1
      when "001001101000" =>  data <= "00000010";  -- 268 = 2
      when "001001101001" =>  data <= "11110000";  -- 269 = F0
      when "001001101010" =>  data <= "00000101";  -- 26A = 5
      when "001001101011" =>  data <= "10101001";  -- 26B = A9
      when "001001101100" =>  data <= "00110001";  -- 26C = 31
      when "001001101101" =>  data <= "01001100";  -- 26D = 4C
      when "001001101110" =>  data <= "01000001";  -- 26E = 41
      when "001001101111" =>  data <= "11111001";  -- 26F = F9
      when "001001110000" =>  data <= "10101001";  -- 270 = A9
      when "001001110001" =>  data <= "10001101";  -- 271 = 8D
      when "001001110010" =>  data <= "10001101";  -- 272 = 8D
      when "001001110011" =>  data <= "00000001";  -- 273 = 1
      when "001001110100" =>  data <= "00000010";  -- 274 = 2
      when "001001110101" =>  data <= "10101001";  -- 275 = A9
      when "001001110110" =>  data <= "10011000";  -- 276 = 98
      when "001001110111" =>  data <= "10001101";  -- 277 = 8D
      when "001001111000" =>  data <= "00000000";  -- 278 = 0
      when "001001111001" =>  data <= "00000010";  -- 279 = 2
      when "001001111010" =>  data <= "10101001";  -- 27A = A9
      when "001001111011" =>  data <= "11110100";  -- 27B = F4
      when "001001111100" =>  data <= "00111000";  -- 27C = 38
      when "001001111101" =>  data <= "01101101";  -- 27D = 6D
      when "001001111110" =>  data <= "00000000";  -- 27E = 0
      when "001001111111" =>  data <= "00000010";  -- 27F = 2
      when "001010000000" =>  data <= "11001101";  -- 280 = CD
      when "001010000001" =>  data <= "00000001";  -- 281 = 1
      when "001010000010" =>  data <= "00000010";  -- 282 = 2
      when "001010000011" =>  data <= "11110000";  -- 283 = F0
      when "001010000100" =>  data <= "00000101";  -- 284 = 5
      when "001010000101" =>  data <= "10101001";  -- 285 = A9
      when "001010000110" =>  data <= "00110010";  -- 286 = 32
      when "001010000111" =>  data <= "01001100";  -- 287 = 4C
      when "001010001000" =>  data <= "01000001";  -- 288 = 41
      when "001010001001" =>  data <= "11111001";  -- 289 = F9
      when "001010001010" =>  data <= "10101001";  -- 28A = A9
      when "001010001011" =>  data <= "00100011";  -- 28B = 23
      when "001010001100" =>  data <= "10001101";  -- 28C = 8D
      when "001010001101" =>  data <= "00000001";  -- 28D = 1
      when "001010001110" =>  data <= "10000000";  -- 28E = 80
      when "001010001111" =>  data <= "10100000";  -- 28F = A0
      when "001010010000" =>  data <= "10000100";  -- 290 = 84
      when "001010010001" =>  data <= "10001100";  -- 291 = 8C
      when "001010010010" =>  data <= "00000001";  -- 292 = 1
      when "001010010011" =>  data <= "00000010";  -- 293 = 2
      when "001010010100" =>  data <= "10100010";  -- 294 = A2
      when "001010010101" =>  data <= "10110100";  -- 295 = B4
      when "001010010110" =>  data <= "10001110";  -- 296 = 8E
      when "001010010111" =>  data <= "00000000";  -- 297 = 0
      when "001010011000" =>  data <= "00000010";  -- 298 = 2
      when "001010011001" =>  data <= "10101001";  -- 299 = A9
      when "001010011010" =>  data <= "10000110";  -- 29A = 86
      when "001010011011" =>  data <= "00101101";  -- 29B = 2D
      when "001010011100" =>  data <= "00000000";  -- 29C = 0
      when "001010011101" =>  data <= "00000010";  -- 29D = 2
      when "001010011110" =>  data <= "11001101";  -- 29E = CD
      when "001010011111" =>  data <= "00000001";  -- 29F = 1
      when "001010100000" =>  data <= "00000010";  -- 2A0 = 2
      when "001010100001" =>  data <= "11110000";  -- 2A1 = F0
      when "001010100010" =>  data <= "00000101";  -- 2A2 = 5
      when "001010100011" =>  data <= "10101001";  -- 2A3 = A9
      when "001010100100" =>  data <= "00110011";  -- 2A4 = 33
      when "001010100101" =>  data <= "01001100";  -- 2A5 = 4C
      when "001010100110" =>  data <= "01000001";  -- 2A6 = 41
      when "001010100111" =>  data <= "11111001";  -- 2A7 = F9
      when "001010101000" =>  data <= "10101001";  -- 2A8 = A9
      when "001010101001" =>  data <= "00100100";  -- 2A9 = 24
      when "001010101010" =>  data <= "10001101";  -- 2AA = 8D
      when "001010101011" =>  data <= "00000001";  -- 2AB = 1
      when "001010101100" =>  data <= "10000000";  -- 2AC = 80
      when "001010101101" =>  data <= "10100010";  -- 2AD = A2
      when "001010101110" =>  data <= "01010101";  -- 2AE = 55
      when "001010101111" =>  data <= "10001110";  -- 2AF = 8E
      when "001010110000" =>  data <= "00000000";  -- 2B0 = 0
      when "001010110001" =>  data <= "00000010";  -- 2B1 = 2
      when "001010110010" =>  data <= "00001110";  -- 2B2 = E
      when "001010110011" =>  data <= "00000000";  -- 2B3 = 0
      when "001010110100" =>  data <= "00000010";  -- 2B4 = 2
      when "001010110101" =>  data <= "10101101";  -- 2B5 = AD
      when "001010110110" =>  data <= "00000000";  -- 2B6 = 0
      when "001010110111" =>  data <= "00000010";  -- 2B7 = 2
      when "001010111000" =>  data <= "11001001";  -- 2B8 = C9
      when "001010111001" =>  data <= "10101010";  -- 2B9 = AA
      when "001010111010" =>  data <= "11110000";  -- 2BA = F0
      when "001010111011" =>  data <= "00000101";  -- 2BB = 5
      when "001010111100" =>  data <= "10101001";  -- 2BC = A9
      when "001010111101" =>  data <= "00110100";  -- 2BD = 34
      when "001010111110" =>  data <= "01001100";  -- 2BE = 4C
      when "001010111111" =>  data <= "01000001";  -- 2BF = 41
      when "001011000000" =>  data <= "11111001";  -- 2C0 = F9
      when "001011000001" =>  data <= "10101001";  -- 2C1 = A9
      when "001011000010" =>  data <= "00100101";  -- 2C2 = 25
      when "001011000011" =>  data <= "10001101";  -- 2C3 = 8D
      when "001011000100" =>  data <= "00000001";  -- 2C4 = 1
      when "001011000101" =>  data <= "10000000";  -- 2C5 = 80
      when "001011000110" =>  data <= "10101001";  -- 2C6 = A9
      when "001011000111" =>  data <= "01010011";  -- 2C7 = 53
      when "001011001000" =>  data <= "10001101";  -- 2C8 = 8D
      when "001011001001" =>  data <= "00000000";  -- 2C9 = 0
      when "001011001010" =>  data <= "00000010";  -- 2CA = 2
      when "001011001011" =>  data <= "10101001";  -- 2CB = A9
      when "001011001100" =>  data <= "00000000";  -- 2CC = 0
      when "001011001101" =>  data <= "10100010";  -- 2CD = A2
      when "001011001110" =>  data <= "01010011";  -- 2CE = 53
      when "001011001111" =>  data <= "11101100";  -- 2CF = EC
      when "001011010000" =>  data <= "00000000";  -- 2D0 = 0
      when "001011010001" =>  data <= "00000010";  -- 2D1 = 2
      when "001011010010" =>  data <= "11110000";  -- 2D2 = F0
      when "001011010011" =>  data <= "00000101";  -- 2D3 = 5
      when "001011010100" =>  data <= "10101001";  -- 2D4 = A9
      when "001011010101" =>  data <= "00110101";  -- 2D5 = 35
      when "001011010110" =>  data <= "01001100";  -- 2D6 = 4C
      when "001011010111" =>  data <= "01000001";  -- 2D7 = 41
      when "001011011000" =>  data <= "11111001";  -- 2D8 = F9
      when "001011011001" =>  data <= "10101001";  -- 2D9 = A9
      when "001011011010" =>  data <= "00100110";  -- 2DA = 26
      when "001011011011" =>  data <= "10001101";  -- 2DB = 8D
      when "001011011100" =>  data <= "00000001";  -- 2DC = 1
      when "001011011101" =>  data <= "10000000";  -- 2DD = 80
      when "001011011110" =>  data <= "10101001";  -- 2DE = A9
      when "001011011111" =>  data <= "01000101";  -- 2DF = 45
      when "001011100000" =>  data <= "10001101";  -- 2E0 = 8D
      when "001011100001" =>  data <= "00000000";  -- 2E1 = 0
      when "001011100010" =>  data <= "00000010";  -- 2E2 = 2
      when "001011100011" =>  data <= "10101001";  -- 2E3 = A9
      when "001011100100" =>  data <= "00000000";  -- 2E4 = 0
      when "001011100101" =>  data <= "10100000";  -- 2E5 = A0
      when "001011100110" =>  data <= "01000101";  -- 2E6 = 45
      when "001011100111" =>  data <= "11001100";  -- 2E7 = CC
      when "001011101000" =>  data <= "00000000";  -- 2E8 = 0
      when "001011101001" =>  data <= "00000010";  -- 2E9 = 2
      when "001011101010" =>  data <= "11110000";  -- 2EA = F0
      when "001011101011" =>  data <= "00000101";  -- 2EB = 5
      when "001011101100" =>  data <= "10101001";  -- 2EC = A9
      when "001011101101" =>  data <= "00110110";  -- 2ED = 36
      when "001011101110" =>  data <= "01001100";  -- 2EE = 4C
      when "001011101111" =>  data <= "01000001";  -- 2EF = 41
      when "001011110000" =>  data <= "11111001";  -- 2F0 = F9
      when "001011110001" =>  data <= "10101001";  -- 2F1 = A9
      when "001011110010" =>  data <= "00100111";  -- 2F2 = 27
      when "001011110011" =>  data <= "10001101";  -- 2F3 = 8D
      when "001011110100" =>  data <= "00000001";  -- 2F4 = 1
      when "001011110101" =>  data <= "10000000";  -- 2F5 = 80
      when "001011110110" =>  data <= "10101001";  -- 2F6 = A9
      when "001011110111" =>  data <= "11101111";  -- 2F7 = EF
      when "001011111000" =>  data <= "10001101";  -- 2F8 = 8D
      when "001011111001" =>  data <= "00000000";  -- 2F9 = 0
      when "001011111010" =>  data <= "00000010";  -- 2FA = 2
      when "001011111011" =>  data <= "11001110";  -- 2FB = CE
      when "001011111100" =>  data <= "00000000";  -- 2FC = 0
      when "001011111101" =>  data <= "00000010";  -- 2FD = 2
      when "001011111110" =>  data <= "10101001";  -- 2FE = A9
      when "001011111111" =>  data <= "11101110";  -- 2FF = EE
      when "001100000000" =>  data <= "11001101";  -- 300 = CD
      when "001100000001" =>  data <= "00000000";  -- 301 = 0
      when "001100000010" =>  data <= "00000010";  -- 302 = 2
      when "001100000011" =>  data <= "11110000";  -- 303 = F0
      when "001100000100" =>  data <= "00000101";  -- 304 = 5
      when "001100000101" =>  data <= "10101001";  -- 305 = A9
      when "001100000110" =>  data <= "00110111";  -- 306 = 37
      when "001100000111" =>  data <= "01001100";  -- 307 = 4C
      when "001100001000" =>  data <= "01000001";  -- 308 = 41
      when "001100001001" =>  data <= "11111001";  -- 309 = F9
      when "001100001010" =>  data <= "10101001";  -- 30A = A9
      when "001100001011" =>  data <= "00000001";  -- 30B = 1
      when "001100001100" =>  data <= "10001101";  -- 30C = 8D
      when "001100001101" =>  data <= "00000000";  -- 30D = 0
      when "001100001110" =>  data <= "00000010";  -- 30E = 2
      when "001100001111" =>  data <= "11001110";  -- 30F = CE
      when "001100010000" =>  data <= "00000000";  -- 310 = 0
      when "001100010001" =>  data <= "00000010";  -- 311 = 2
      when "001100010010" =>  data <= "11110000";  -- 312 = F0
      when "001100010011" =>  data <= "00000101";  -- 313 = 5
      when "001100010100" =>  data <= "10101001";  -- 314 = A9
      when "001100010101" =>  data <= "00111000";  -- 315 = 38
      when "001100010110" =>  data <= "01001100";  -- 316 = 4C
      when "001100010111" =>  data <= "01000001";  -- 317 = 41
      when "001100011000" =>  data <= "11111001";  -- 318 = F9
      when "001100011001" =>  data <= "10101001";  -- 319 = A9
      when "001100011010" =>  data <= "00101000";  -- 31A = 28
      when "001100011011" =>  data <= "10001101";  -- 31B = 8D
      when "001100011100" =>  data <= "00000001";  -- 31C = 1
      when "001100011101" =>  data <= "10000000";  -- 31D = 80
      when "001100011110" =>  data <= "10101001";  -- 31E = A9
      when "001100011111" =>  data <= "11101111";  -- 31F = EF
      when "001100100000" =>  data <= "10001101";  -- 320 = 8D
      when "001100100001" =>  data <= "00000000";  -- 321 = 0
      when "001100100010" =>  data <= "00000010";  -- 322 = 2
      when "001100100011" =>  data <= "11101110";  -- 323 = EE
      when "001100100100" =>  data <= "00000000";  -- 324 = 0
      when "001100100101" =>  data <= "00000010";  -- 325 = 2
      when "001100100110" =>  data <= "10101001";  -- 326 = A9
      when "001100100111" =>  data <= "11110000";  -- 327 = F0
      when "001100101000" =>  data <= "11001101";  -- 328 = CD
      when "001100101001" =>  data <= "00000000";  -- 329 = 0
      when "001100101010" =>  data <= "00000010";  -- 32A = 2
      when "001100101011" =>  data <= "11110000";  -- 32B = F0
      when "001100101100" =>  data <= "00000101";  -- 32C = 5
      when "001100101101" =>  data <= "10101001";  -- 32D = A9
      when "001100101110" =>  data <= "00111001";  -- 32E = 39
      when "001100101111" =>  data <= "01001100";  -- 32F = 4C
      when "001100110000" =>  data <= "01000001";  -- 330 = 41
      when "001100110001" =>  data <= "11111001";  -- 331 = F9
      when "001100110010" =>  data <= "10101001";  -- 332 = A9
      when "001100110011" =>  data <= "11111111";  -- 333 = FF
      when "001100110100" =>  data <= "10001101";  -- 334 = 8D
      when "001100110101" =>  data <= "00000000";  -- 335 = 0
      when "001100110110" =>  data <= "00000010";  -- 336 = 2
      when "001100110111" =>  data <= "11101110";  -- 337 = EE
      when "001100111000" =>  data <= "00000000";  -- 338 = 0
      when "001100111001" =>  data <= "00000010";  -- 339 = 2
      when "001100111010" =>  data <= "11110000";  -- 33A = F0
      when "001100111011" =>  data <= "00000101";  -- 33B = 5
      when "001100111100" =>  data <= "10101001";  -- 33C = A9
      when "001100111101" =>  data <= "01000000";  -- 33D = 40
      when "001100111110" =>  data <= "01001100";  -- 33E = 4C
      when "001100111111" =>  data <= "01000001";  -- 33F = 41
      when "001101000000" =>  data <= "11111001";  -- 340 = F9
      when "001101000001" =>  data <= "10101001";  -- 341 = A9
      when "001101000010" =>  data <= "00101001";  -- 342 = 29
      when "001101000011" =>  data <= "10001101";  -- 343 = 8D
      when "001101000100" =>  data <= "00000001";  -- 344 = 1
      when "001101000101" =>  data <= "10000000";  -- 345 = 80
      when "001101000110" =>  data <= "10100000";  -- 346 = A0
      when "001101000111" =>  data <= "00110010";  -- 347 = 32
      when "001101001000" =>  data <= "10001100";  -- 348 = 8C
      when "001101001001" =>  data <= "00000001";  -- 349 = 1
      when "001101001010" =>  data <= "00000010";  -- 34A = 2
      when "001101001011" =>  data <= "10100010";  -- 34B = A2
      when "001101001100" =>  data <= "10110100";  -- 34C = B4
      when "001101001101" =>  data <= "10001110";  -- 34D = 8E
      when "001101001110" =>  data <= "00000000";  -- 34E = 0
      when "001101001111" =>  data <= "00000010";  -- 34F = 2
      when "001101010000" =>  data <= "10101001";  -- 350 = A9
      when "001101010001" =>  data <= "10000110";  -- 351 = 86
      when "001101010010" =>  data <= "01001101";  -- 352 = 4D
      when "001101010011" =>  data <= "00000000";  -- 353 = 0
      when "001101010100" =>  data <= "00000010";  -- 354 = 2
      when "001101010101" =>  data <= "11001101";  -- 355 = CD
      when "001101010110" =>  data <= "00000001";  -- 356 = 1
      when "001101010111" =>  data <= "00000010";  -- 357 = 2
      when "001101011000" =>  data <= "11110000";  -- 358 = F0
      when "001101011001" =>  data <= "00000101";  -- 359 = 5
      when "001101011010" =>  data <= "10101001";  -- 35A = A9
      when "001101011011" =>  data <= "01000001";  -- 35B = 41
      when "001101011100" =>  data <= "01001100";  -- 35C = 4C
      when "001101011101" =>  data <= "01000001";  -- 35D = 41
      when "001101011110" =>  data <= "11111001";  -- 35E = F9
      when "001101011111" =>  data <= "10101001";  -- 35F = A9
      when "001101100000" =>  data <= "00101010";  -- 360 = 2A
      when "001101100001" =>  data <= "10001101";  -- 361 = 8D
      when "001101100010" =>  data <= "00000001";  -- 362 = 1
      when "001101100011" =>  data <= "10000000";  -- 363 = 80
      when "001101100100" =>  data <= "10100000";  -- 364 = A0
      when "001101100101" =>  data <= "10110110";  -- 365 = B6
      when "001101100110" =>  data <= "10001100";  -- 366 = 8C
      when "001101100111" =>  data <= "00000001";  -- 367 = 1
      when "001101101000" =>  data <= "00000010";  -- 368 = 2
      when "001101101001" =>  data <= "10100010";  -- 369 = A2
      when "001101101010" =>  data <= "10110100";  -- 36A = B4
      when "001101101011" =>  data <= "10001110";  -- 36B = 8E
      when "001101101100" =>  data <= "00000000";  -- 36C = 0
      when "001101101101" =>  data <= "00000010";  -- 36D = 2
      when "001101101110" =>  data <= "10101001";  -- 36E = A9
      when "001101101111" =>  data <= "10000110";  -- 36F = 86
      when "001101110000" =>  data <= "00001101";  -- 370 = D
      when "001101110001" =>  data <= "00000000";  -- 371 = 0
      when "001101110010" =>  data <= "00000010";  -- 372 = 2
      when "001101110011" =>  data <= "11001101";  -- 373 = CD
      when "001101110100" =>  data <= "00000001";  -- 374 = 1
      when "001101110101" =>  data <= "00000010";  -- 375 = 2
      when "001101110110" =>  data <= "11110000";  -- 376 = F0
      when "001101110111" =>  data <= "00000101";  -- 377 = 5
      when "001101111000" =>  data <= "10101001";  -- 378 = A9
      when "001101111001" =>  data <= "01000010";  -- 379 = 42
      when "001101111010" =>  data <= "01001100";  -- 37A = 4C
      when "001101111011" =>  data <= "01000001";  -- 37B = 41
      when "001101111100" =>  data <= "11111001";  -- 37C = F9
      when "001101111101" =>  data <= "10101001";  -- 37D = A9
      when "001101111110" =>  data <= "00101011";  -- 37E = 2B
      when "001101111111" =>  data <= "10001101";  -- 37F = 8D
      when "001110000000" =>  data <= "00000001";  -- 380 = 1
      when "001110000001" =>  data <= "10000000";  -- 381 = 80
      when "001110000010" =>  data <= "00011000";  -- 382 = 18
      when "001110000011" =>  data <= "10100010";  -- 383 = A2
      when "001110000100" =>  data <= "10101010";  -- 384 = AA
      when "001110000101" =>  data <= "10001110";  -- 385 = 8E
      when "001110000110" =>  data <= "00000000";  -- 386 = 0
      when "001110000111" =>  data <= "00000010";  -- 387 = 2
      when "001110001000" =>  data <= "00101110";  -- 388 = 2E
      when "001110001001" =>  data <= "00000000";  -- 389 = 0
      when "001110001010" =>  data <= "00000010";  -- 38A = 2
      when "001110001011" =>  data <= "10110000";  -- 38B = B0
      when "001110001100" =>  data <= "00000101";  -- 38C = 5
      when "001110001101" =>  data <= "10101001";  -- 38D = A9
      when "001110001110" =>  data <= "01000011";  -- 38E = 43
      when "001110001111" =>  data <= "01001100";  -- 38F = 4C
      when "001110010000" =>  data <= "01000001";  -- 390 = 41
      when "001110010001" =>  data <= "11111001";  -- 391 = F9
      when "001110010010" =>  data <= "10101101";  -- 392 = AD
      when "001110010011" =>  data <= "00000000";  -- 393 = 0
      when "001110010100" =>  data <= "00000010";  -- 394 = 2
      when "001110010101" =>  data <= "11001001";  -- 395 = C9
      when "001110010110" =>  data <= "01010100";  -- 396 = 54
      when "001110010111" =>  data <= "11110000";  -- 397 = F0
      when "001110011000" =>  data <= "00000101";  -- 398 = 5
      when "001110011001" =>  data <= "10101001";  -- 399 = A9
      when "001110011010" =>  data <= "01000100";  -- 39A = 44
      when "001110011011" =>  data <= "01001100";  -- 39B = 4C
      when "001110011100" =>  data <= "01000001";  -- 39C = 41
      when "001110011101" =>  data <= "11111001";  -- 39D = F9
      when "001110011110" =>  data <= "10101001";  -- 39E = A9
      when "001110011111" =>  data <= "00101100";  -- 39F = 2C
      when "001110100000" =>  data <= "10001101";  -- 3A0 = 8D
      when "001110100001" =>  data <= "00000001";  -- 3A1 = 1
      when "001110100010" =>  data <= "10000000";  -- 3A2 = 80
      when "001110100011" =>  data <= "00011000";  -- 3A3 = 18
      when "001110100100" =>  data <= "10100010";  -- 3A4 = A2
      when "001110100101" =>  data <= "01010101";  -- 3A5 = 55
      when "001110100110" =>  data <= "10001110";  -- 3A6 = 8E
      when "001110100111" =>  data <= "00000000";  -- 3A7 = 0
      when "001110101000" =>  data <= "00000010";  -- 3A8 = 2
      when "001110101001" =>  data <= "01101110";  -- 3A9 = 6E
      when "001110101010" =>  data <= "00000000";  -- 3AA = 0
      when "001110101011" =>  data <= "00000010";  -- 3AB = 2
      when "001110101100" =>  data <= "10110000";  -- 3AC = B0
      when "001110101101" =>  data <= "00000101";  -- 3AD = 5
      when "001110101110" =>  data <= "10101001";  -- 3AE = A9
      when "001110101111" =>  data <= "01000101";  -- 3AF = 45
      when "001110110000" =>  data <= "01001100";  -- 3B0 = 4C
      when "001110110001" =>  data <= "01000001";  -- 3B1 = 41
      when "001110110010" =>  data <= "11111001";  -- 3B2 = F9
      when "001110110011" =>  data <= "10101101";  -- 3B3 = AD
      when "001110110100" =>  data <= "00000000";  -- 3B4 = 0
      when "001110110101" =>  data <= "00000010";  -- 3B5 = 2
      when "001110110110" =>  data <= "11001001";  -- 3B6 = C9
      when "001110110111" =>  data <= "00101010";  -- 3B7 = 2A
      when "001110111000" =>  data <= "11110000";  -- 3B8 = F0
      when "001110111001" =>  data <= "00000101";  -- 3B9 = 5
      when "001110111010" =>  data <= "10101001";  -- 3BA = A9
      when "001110111011" =>  data <= "01000110";  -- 3BB = 46
      when "001110111100" =>  data <= "01001100";  -- 3BC = 4C
      when "001110111101" =>  data <= "01000001";  -- 3BD = 41
      when "001110111110" =>  data <= "11111001";  -- 3BE = F9
      when "001110111111" =>  data <= "10101001";  -- 3BF = A9
      when "001111000000" =>  data <= "00101101";  -- 3C0 = 2D
      when "001111000001" =>  data <= "10001101";  -- 3C1 = 8D
      when "001111000010" =>  data <= "00000001";  -- 3C2 = 1
      when "001111000011" =>  data <= "10000000";  -- 3C3 = 80
      when "001111000100" =>  data <= "10100010";  -- 3C4 = A2
      when "001111000101" =>  data <= "10010110";  -- 3C5 = 96
      when "001111000110" =>  data <= "10001110";  -- 3C6 = 8E
      when "001111000111" =>  data <= "00000000";  -- 3C7 = 0
      when "001111001000" =>  data <= "00000010";  -- 3C8 = 2
      when "001111001001" =>  data <= "01001110";  -- 3C9 = 4E
      when "001111001010" =>  data <= "00000000";  -- 3CA = 0
      when "001111001011" =>  data <= "00000010";  -- 3CB = 2
      when "001111001100" =>  data <= "10101101";  -- 3CC = AD
      when "001111001101" =>  data <= "00000000";  -- 3CD = 0
      when "001111001110" =>  data <= "00000010";  -- 3CE = 2
      when "001111001111" =>  data <= "11001001";  -- 3CF = C9
      when "001111010000" =>  data <= "01001011";  -- 3D0 = 4B
      when "001111010001" =>  data <= "11110000";  -- 3D1 = F0
      when "001111010010" =>  data <= "00000101";  -- 3D2 = 5
      when "001111010011" =>  data <= "10101001";  -- 3D3 = A9
      when "001111010100" =>  data <= "01000111";  -- 3D4 = 47
      when "001111010101" =>  data <= "01001100";  -- 3D5 = 4C
      when "001111010110" =>  data <= "01000001";  -- 3D6 = 41
      when "001111010111" =>  data <= "11111001";  -- 3D7 = F9
      when "001111011000" =>  data <= "10101001";  -- 3D8 = A9
      when "001111011001" =>  data <= "00101110";  -- 3D9 = 2E
      when "001111011010" =>  data <= "10001101";  -- 3DA = 8D
      when "001111011011" =>  data <= "00000001";  -- 3DB = 1
      when "001111011100" =>  data <= "10000000";  -- 3DC = 80
      when "001111011101" =>  data <= "10100010";  -- 3DD = A2
      when "001111011110" =>  data <= "01000010";  -- 3DE = 42
      when "001111011111" =>  data <= "10001110";  -- 3DF = 8E
      when "001111100000" =>  data <= "00000000";  -- 3E0 = 0
      when "001111100001" =>  data <= "00000010";  -- 3E1 = 2
      when "001111100010" =>  data <= "10100010";  -- 3E2 = A2
      when "001111100011" =>  data <= "10011111";  -- 3E3 = 9F
      when "001111100100" =>  data <= "10001110";  -- 3E4 = 8E
      when "001111100101" =>  data <= "00000001";  -- 3E5 = 1
      when "001111100110" =>  data <= "00000010";  -- 3E6 = 2
      when "001111100111" =>  data <= "10101110";  -- 3E7 = AE
      when "001111101000" =>  data <= "00000000";  -- 3E8 = 0
      when "001111101001" =>  data <= "00000010";  -- 3E9 = 2
      when "001111101010" =>  data <= "11100000";  -- 3EA = E0
      when "001111101011" =>  data <= "01000010";  -- 3EB = 42
      when "001111101100" =>  data <= "11110000";  -- 3EC = F0
      when "001111101101" =>  data <= "00000101";  -- 3ED = 5
      when "001111101110" =>  data <= "10101001";  -- 3EE = A9
      when "001111101111" =>  data <= "01001000";  -- 3EF = 48
      when "001111110000" =>  data <= "01001100";  -- 3F0 = 4C
      when "001111110001" =>  data <= "01000001";  -- 3F1 = 41
      when "001111110010" =>  data <= "11111001";  -- 3F2 = F9
      when "001111110011" =>  data <= "10101110";  -- 3F3 = AE
      when "001111110100" =>  data <= "00000001";  -- 3F4 = 1
      when "001111110101" =>  data <= "00000010";  -- 3F5 = 2
      when "001111110110" =>  data <= "11100000";  -- 3F6 = E0
      when "001111110111" =>  data <= "10011111";  -- 3F7 = 9F
      when "001111111000" =>  data <= "11110000";  -- 3F8 = F0
      when "001111111001" =>  data <= "00000101";  -- 3F9 = 5
      when "001111111010" =>  data <= "10101001";  -- 3FA = A9
      when "001111111011" =>  data <= "01001001";  -- 3FB = 49
      when "001111111100" =>  data <= "01001100";  -- 3FC = 4C
      when "001111111101" =>  data <= "01000001";  -- 3FD = 41
      when "001111111110" =>  data <= "11111001";  -- 3FE = F9
      when "001111111111" =>  data <= "10101001";  -- 3FF = A9
      when "010000000000" =>  data <= "00101111";  -- 400 = 2F
      when "010000000001" =>  data <= "10001101";  -- 401 = 8D
      when "010000000010" =>  data <= "00000001";  -- 402 = 1
      when "010000000011" =>  data <= "10000000";  -- 403 = 80
      when "010000000100" =>  data <= "10100000";  -- 404 = A0
      when "010000000101" =>  data <= "00110100";  -- 405 = 34
      when "010000000110" =>  data <= "10001100";  -- 406 = 8C
      when "010000000111" =>  data <= "00000000";  -- 407 = 0
      when "010000001000" =>  data <= "00000010";  -- 408 = 2
      when "010000001001" =>  data <= "10100000";  -- 409 = A0
      when "010000001010" =>  data <= "01110101";  -- 40A = 75
      when "010000001011" =>  data <= "10001100";  -- 40B = 8C
      when "010000001100" =>  data <= "00000001";  -- 40C = 1
      when "010000001101" =>  data <= "00000010";  -- 40D = 2
      when "010000001110" =>  data <= "10101100";  -- 40E = AC
      when "010000001111" =>  data <= "00000000";  -- 40F = 0
      when "010000010000" =>  data <= "00000010";  -- 410 = 2
      when "010000010001" =>  data <= "11000000";  -- 411 = C0
      when "010000010010" =>  data <= "00110100";  -- 412 = 34
      when "010000010011" =>  data <= "11110000";  -- 413 = F0
      when "010000010100" =>  data <= "00000101";  -- 414 = 5
      when "010000010101" =>  data <= "10101001";  -- 415 = A9
      when "010000010110" =>  data <= "01001010";  -- 416 = 4A
      when "010000010111" =>  data <= "01001100";  -- 417 = 4C
      when "010000011000" =>  data <= "01000001";  -- 418 = 41
      when "010000011001" =>  data <= "11111001";  -- 419 = F9
      when "010000011010" =>  data <= "10101100";  -- 41A = AC
      when "010000011011" =>  data <= "00000001";  -- 41B = 1
      when "010000011100" =>  data <= "00000010";  -- 41C = 2
      when "010000011101" =>  data <= "11000000";  -- 41D = C0
      when "010000011110" =>  data <= "01110101";  -- 41E = 75
      when "010000011111" =>  data <= "11110000";  -- 41F = F0
      when "010000100000" =>  data <= "00000101";  -- 420 = 5
      when "010000100001" =>  data <= "10101001";  -- 421 = A9
      when "010000100010" =>  data <= "01001011";  -- 422 = 4B
      when "010000100011" =>  data <= "01001100";  -- 423 = 4C
      when "010000100100" =>  data <= "01000001";  -- 424 = 41
      when "010000100101" =>  data <= "11111001";  -- 425 = F9
      when "010000100110" =>  data <= "10101001";  -- 426 = A9
      when "010000100111" =>  data <= "00110000";  -- 427 = 30
      when "010000101000" =>  data <= "10001101";  -- 428 = 8D
      when "010000101001" =>  data <= "00000001";  -- 429 = 1
      when "010000101010" =>  data <= "10000000";  -- 42A = 80
      when "010000101011" =>  data <= "10101001";  -- 42B = A9
      when "010000101100" =>  data <= "00010010";  -- 42C = 12
      when "010000101101" =>  data <= "10001101";  -- 42D = 8D
      when "010000101110" =>  data <= "00000001";  -- 42E = 1
      when "010000101111" =>  data <= "00000010";  -- 42F = 2
      when "010000110000" =>  data <= "10101001";  -- 430 = A9
      when "010000110001" =>  data <= "01000001";  -- 431 = 41
      when "010000110010" =>  data <= "10001101";  -- 432 = 8D
      when "010000110011" =>  data <= "00000000";  -- 433 = 0
      when "010000110100" =>  data <= "00000010";  -- 434 = 2
      when "010000110101" =>  data <= "10101001";  -- 435 = A9
      when "010000110110" =>  data <= "01010011";  -- 436 = 53
      when "010000110111" =>  data <= "00111000";  -- 437 = 38
      when "010000111000" =>  data <= "11101101";  -- 438 = ED
      when "010000111001" =>  data <= "00000000";  -- 439 = 0
      when "010000111010" =>  data <= "00000010";  -- 43A = 2
      when "010000111011" =>  data <= "11001101";  -- 43B = CD
      when "010000111100" =>  data <= "00000001";  -- 43C = 1
      when "010000111101" =>  data <= "00000010";  -- 43D = 2
      when "010000111110" =>  data <= "11110000";  -- 43E = F0
      when "010000111111" =>  data <= "00000101";  -- 43F = 5
      when "010001000000" =>  data <= "10101001";  -- 440 = A9
      when "010001000001" =>  data <= "01001100";  -- 441 = 4C
      when "010001000010" =>  data <= "01001100";  -- 442 = 4C
      when "010001000011" =>  data <= "01000001";  -- 443 = 41
      when "010001000100" =>  data <= "11111001";  -- 444 = F9
      when "010001000101" =>  data <= "10101001";  -- 445 = A9
      when "010001000110" =>  data <= "01011011";  -- 446 = 5B
      when "010001000111" =>  data <= "10001101";  -- 447 = 8D
      when "010001001000" =>  data <= "00000001";  -- 448 = 1
      when "010001001001" =>  data <= "00000010";  -- 449 = 2
      when "010001001010" =>  data <= "10101001";  -- 44A = A9
      when "010001001011" =>  data <= "10011000";  -- 44B = 98
      when "010001001100" =>  data <= "10001101";  -- 44C = 8D
      when "010001001101" =>  data <= "00000000";  -- 44D = 0
      when "010001001110" =>  data <= "00000010";  -- 44E = 2
      when "010001001111" =>  data <= "10101001";  -- 44F = A9
      when "010001010000" =>  data <= "11110100";  -- 450 = F4
      when "010001010001" =>  data <= "00011000";  -- 451 = 18
      when "010001010010" =>  data <= "11101101";  -- 452 = ED
      when "010001010011" =>  data <= "00000000";  -- 453 = 0
      when "010001010100" =>  data <= "00000010";  -- 454 = 2
      when "010001010101" =>  data <= "11001101";  -- 455 = CD
      when "010001010110" =>  data <= "00000001";  -- 456 = 1
      when "010001010111" =>  data <= "00000010";  -- 457 = 2
      when "010001011000" =>  data <= "11110000";  -- 458 = F0
      when "010001011001" =>  data <= "00000101";  -- 459 = 5
      when "010001011010" =>  data <= "10101001";  -- 45A = A9
      when "010001011011" =>  data <= "01001101";  -- 45B = 4D
      when "010001011100" =>  data <= "01001100";  -- 45C = 4C
      when "010001011101" =>  data <= "01000001";  -- 45D = 41
      when "010001011110" =>  data <= "11111001";  -- 45E = F9
      when "010001011111" =>  data <= "10101001";  -- 45F = A9
      when "010001100000" =>  data <= "00110001";  -- 460 = 31
      when "010001100001" =>  data <= "10001101";  -- 461 = 8D
      when "010001100010" =>  data <= "00000001";  -- 462 = 1
      when "010001100011" =>  data <= "10000000";  -- 463 = 80
      when "010001100100" =>  data <= "10101001";  -- 464 = A9
      when "010001100101" =>  data <= "01000010";  -- 465 = 42
      when "010001100110" =>  data <= "01001000";  -- 466 = 48
      when "010001100111" =>  data <= "10101001";  -- 467 = A9
      when "010001101000" =>  data <= "11101101";  -- 468 = ED
      when "010001101001" =>  data <= "01001000";  -- 469 = 48
      when "010001101010" =>  data <= "10101001";  -- 46A = A9
      when "010001101011" =>  data <= "10111110";  -- 46B = BE
      when "010001101100" =>  data <= "01001000";  -- 46C = 48
      when "010001101101" =>  data <= "10101001";  -- 46D = A9
      when "010001101110" =>  data <= "00000000";  -- 46E = 0
      when "010001101111" =>  data <= "01101000";  -- 46F = 68
      when "010001110000" =>  data <= "11001001";  -- 470 = C9
      when "010001110001" =>  data <= "10111110";  -- 471 = BE
      when "010001110010" =>  data <= "11010000";  -- 472 = D0
      when "010001110011" =>  data <= "00001101";  -- 473 = D
      when "010001110100" =>  data <= "01101000";  -- 474 = 68
      when "010001110101" =>  data <= "11001001";  -- 475 = C9
      when "010001110110" =>  data <= "11101101";  -- 476 = ED
      when "010001110111" =>  data <= "11010000";  -- 477 = D0
      when "010001111000" =>  data <= "00001000";  -- 478 = 8
      when "010001111001" =>  data <= "01101000";  -- 479 = 68
      when "010001111010" =>  data <= "11001001";  -- 47A = C9
      when "010001111011" =>  data <= "01000010";  -- 47B = 42
      when "010001111100" =>  data <= "11010000";  -- 47C = D0
      when "010001111101" =>  data <= "00000011";  -- 47D = 3
      when "010001111110" =>  data <= "01001100";  -- 47E = 4C
      when "010001111111" =>  data <= "10000110";  -- 47F = 86
      when "010010000000" =>  data <= "11110100";  -- 480 = F4
      when "010010000001" =>  data <= "10101001";  -- 481 = A9
      when "010010000010" =>  data <= "01001110";  -- 482 = 4E
      when "010010000011" =>  data <= "01001100";  -- 483 = 4C
      when "010010000100" =>  data <= "01000001";  -- 484 = 41
      when "010010000101" =>  data <= "11111001";  -- 485 = F9
      when "010010000110" =>  data <= "10101001";  -- 486 = A9
      when "010010000111" =>  data <= "00110010";  -- 487 = 32
      when "010010001000" =>  data <= "10001101";  -- 488 = 8D
      when "010010001001" =>  data <= "00000001";  -- 489 = 1
      when "010010001010" =>  data <= "10000000";  -- 48A = 80
      when "010010001011" =>  data <= "10100010";  -- 48B = A2
      when "010010001100" =>  data <= "00000000";  -- 48C = 0
      when "010010001101" =>  data <= "00011000";  -- 48D = 18
      when "010010001110" =>  data <= "10101001";  -- 48E = A9
      when "010010001111" =>  data <= "00000011";  -- 48F = 3
      when "010010010000" =>  data <= "10011101";  -- 490 = 9D
      when "010010010001" =>  data <= "00000000";  -- 491 = 0
      when "010010010010" =>  data <= "00000010";  -- 492 = 2
      when "010010010011" =>  data <= "01101001";  -- 493 = 69
      when "010010010100" =>  data <= "00000111";  -- 494 = 7
      when "010010010101" =>  data <= "11101000";  -- 495 = E8
      when "010010010110" =>  data <= "10011101";  -- 496 = 9D
      when "010010010111" =>  data <= "00000000";  -- 497 = 0
      when "010010011000" =>  data <= "00000010";  -- 498 = 2
      when "010010011001" =>  data <= "01101001";  -- 499 = 69
      when "010010011010" =>  data <= "00000111";  -- 49A = 7
      when "010010011011" =>  data <= "11101000";  -- 49B = E8
      when "010010011100" =>  data <= "10011101";  -- 49C = 9D
      when "010010011101" =>  data <= "00000000";  -- 49D = 0
      when "010010011110" =>  data <= "00000010";  -- 49E = 2
      when "010010011111" =>  data <= "01101001";  -- 49F = 69
      when "010010100000" =>  data <= "00000111";  -- 4A0 = 7
      when "010010100001" =>  data <= "11101000";  -- 4A1 = E8
      when "010010100010" =>  data <= "10011101";  -- 4A2 = 9D
      when "010010100011" =>  data <= "00000000";  -- 4A3 = 0
      when "010010100100" =>  data <= "00000010";  -- 4A4 = 2
      when "010010100101" =>  data <= "01101001";  -- 4A5 = 69
      when "010010100110" =>  data <= "00000111";  -- 4A6 = 7
      when "010010100111" =>  data <= "11101000";  -- 4A7 = E8
      when "010010101000" =>  data <= "10011101";  -- 4A8 = 9D
      when "010010101001" =>  data <= "00000000";  -- 4A9 = 0
      when "010010101010" =>  data <= "00000010";  -- 4AA = 2
      when "010010101011" =>  data <= "01101001";  -- 4AB = 69
      when "010010101100" =>  data <= "00000111";  -- 4AC = 7
      when "010010101101" =>  data <= "11101000";  -- 4AD = E8
      when "010010101110" =>  data <= "10011101";  -- 4AE = 9D
      when "010010101111" =>  data <= "00000000";  -- 4AF = 0
      when "010010110000" =>  data <= "00000010";  -- 4B0 = 2
      when "010010110001" =>  data <= "01101001";  -- 4B1 = 69
      when "010010110010" =>  data <= "00000111";  -- 4B2 = 7
      when "010010110011" =>  data <= "11101000";  -- 4B3 = E8
      when "010010110100" =>  data <= "10011101";  -- 4B4 = 9D
      when "010010110101" =>  data <= "00000000";  -- 4B5 = 0
      when "010010110110" =>  data <= "00000010";  -- 4B6 = 2
      when "010010110111" =>  data <= "10100010";  -- 4B7 = A2
      when "010010111000" =>  data <= "00000000";  -- 4B8 = 0
      when "010010111001" =>  data <= "00011000";  -- 4B9 = 18
      when "010010111010" =>  data <= "10111101";  -- 4BA = BD
      when "010010111011" =>  data <= "00000000";  -- 4BB = 0
      when "010010111100" =>  data <= "00000010";  -- 4BC = 2
      when "010010111101" =>  data <= "11001001";  -- 4BD = C9
      when "010010111110" =>  data <= "00000011";  -- 4BE = 3
      when "010010111111" =>  data <= "11010000";  -- 4BF = D0
      when "010011000000" =>  data <= "00110011";  -- 4C0 = 33
      when "010011000001" =>  data <= "11101000";  -- 4C1 = E8
      when "010011000010" =>  data <= "10111101";  -- 4C2 = BD
      when "010011000011" =>  data <= "00000000";  -- 4C3 = 0
      when "010011000100" =>  data <= "00000010";  -- 4C4 = 2
      when "010011000101" =>  data <= "11001001";  -- 4C5 = C9
      when "010011000110" =>  data <= "00001010";  -- 4C6 = A
      when "010011000111" =>  data <= "11010000";  -- 4C7 = D0
      when "010011001000" =>  data <= "00101011";  -- 4C8 = 2B
      when "010011001001" =>  data <= "11101000";  -- 4C9 = E8
      when "010011001010" =>  data <= "10111101";  -- 4CA = BD
      when "010011001011" =>  data <= "00000000";  -- 4CB = 0
      when "010011001100" =>  data <= "00000010";  -- 4CC = 2
      when "010011001101" =>  data <= "11001001";  -- 4CD = C9
      when "010011001110" =>  data <= "00010001";  -- 4CE = 11
      when "010011001111" =>  data <= "11010000";  -- 4CF = D0
      when "010011010000" =>  data <= "00100011";  -- 4D0 = 23
      when "010011010001" =>  data <= "11101000";  -- 4D1 = E8
      when "010011010010" =>  data <= "10111101";  -- 4D2 = BD
      when "010011010011" =>  data <= "00000000";  -- 4D3 = 0
      when "010011010100" =>  data <= "00000010";  -- 4D4 = 2
      when "010011010101" =>  data <= "11001001";  -- 4D5 = C9
      when "010011010110" =>  data <= "00011000";  -- 4D6 = 18
      when "010011010111" =>  data <= "11010000";  -- 4D7 = D0
      when "010011011000" =>  data <= "00011011";  -- 4D8 = 1B
      when "010011011001" =>  data <= "11101000";  -- 4D9 = E8
      when "010011011010" =>  data <= "10111101";  -- 4DA = BD
      when "010011011011" =>  data <= "00000000";  -- 4DB = 0
      when "010011011100" =>  data <= "00000010";  -- 4DC = 2
      when "010011011101" =>  data <= "11001001";  -- 4DD = C9
      when "010011011110" =>  data <= "00011111";  -- 4DE = 1F
      when "010011011111" =>  data <= "11010000";  -- 4DF = D0
      when "010011100000" =>  data <= "00010011";  -- 4E0 = 13
      when "010011100001" =>  data <= "11101000";  -- 4E1 = E8
      when "010011100010" =>  data <= "10111101";  -- 4E2 = BD
      when "010011100011" =>  data <= "00000000";  -- 4E3 = 0
      when "010011100100" =>  data <= "00000010";  -- 4E4 = 2
      when "010011100101" =>  data <= "11001001";  -- 4E5 = C9
      when "010011100110" =>  data <= "00100110";  -- 4E6 = 26
      when "010011100111" =>  data <= "11010000";  -- 4E7 = D0
      when "010011101000" =>  data <= "00001011";  -- 4E8 = B
      when "010011101001" =>  data <= "11101000";  -- 4E9 = E8
      when "010011101010" =>  data <= "10111101";  -- 4EA = BD
      when "010011101011" =>  data <= "00000000";  -- 4EB = 0
      when "010011101100" =>  data <= "00000010";  -- 4EC = 2
      when "010011101101" =>  data <= "11001001";  -- 4ED = C9
      when "010011101110" =>  data <= "00101101";  -- 4EE = 2D
      when "010011101111" =>  data <= "11010000";  -- 4EF = D0
      when "010011110000" =>  data <= "00000011";  -- 4F0 = 3
      when "010011110001" =>  data <= "01001100";  -- 4F1 = 4C
      when "010011110010" =>  data <= "11111001";  -- 4F2 = F9
      when "010011110011" =>  data <= "11110100";  -- 4F3 = F4
      when "010011110100" =>  data <= "10101001";  -- 4F4 = A9
      when "010011110101" =>  data <= "01001111";  -- 4F5 = 4F
      when "010011110110" =>  data <= "01001100";  -- 4F6 = 4C
      when "010011110111" =>  data <= "01000001";  -- 4F7 = 41
      when "010011111000" =>  data <= "11111001";  -- 4F8 = F9
      when "010011111001" =>  data <= "10101001";  -- 4F9 = A9
      when "010011111010" =>  data <= "00110011";  -- 4FA = 33
      when "010011111011" =>  data <= "10001101";  -- 4FB = 8D
      when "010011111100" =>  data <= "00000001";  -- 4FC = 1
      when "010011111101" =>  data <= "10000000";  -- 4FD = 80
      when "010011111110" =>  data <= "10100000";  -- 4FE = A0
      when "010011111111" =>  data <= "00000000";  -- 4FF = 0
      when "010100000000" =>  data <= "00011000";  -- 500 = 18
      when "010100000001" =>  data <= "10101001";  -- 501 = A9
      when "010100000010" =>  data <= "00000011";  -- 502 = 3
      when "010100000011" =>  data <= "10011001";  -- 503 = 99
      when "010100000100" =>  data <= "00000000";  -- 504 = 0
      when "010100000101" =>  data <= "00000010";  -- 505 = 2
      when "010100000110" =>  data <= "01101001";  -- 506 = 69
      when "010100000111" =>  data <= "00000111";  -- 507 = 7
      when "010100001000" =>  data <= "11001000";  -- 508 = C8
      when "010100001001" =>  data <= "10011001";  -- 509 = 99
      when "010100001010" =>  data <= "00000000";  -- 50A = 0
      when "010100001011" =>  data <= "00000010";  -- 50B = 2
      when "010100001100" =>  data <= "01101001";  -- 50C = 69
      when "010100001101" =>  data <= "00000111";  -- 50D = 7
      when "010100001110" =>  data <= "11001000";  -- 50E = C8
      when "010100001111" =>  data <= "10011001";  -- 50F = 99
      when "010100010000" =>  data <= "00000000";  -- 510 = 0
      when "010100010001" =>  data <= "00000010";  -- 511 = 2
      when "010100010010" =>  data <= "01101001";  -- 512 = 69
      when "010100010011" =>  data <= "00000111";  -- 513 = 7
      when "010100010100" =>  data <= "11001000";  -- 514 = C8
      when "010100010101" =>  data <= "10011001";  -- 515 = 99
      when "010100010110" =>  data <= "00000000";  -- 516 = 0
      when "010100010111" =>  data <= "00000010";  -- 517 = 2
      when "010100011000" =>  data <= "01101001";  -- 518 = 69
      when "010100011001" =>  data <= "00000111";  -- 519 = 7
      when "010100011010" =>  data <= "11001000";  -- 51A = C8
      when "010100011011" =>  data <= "10011001";  -- 51B = 99
      when "010100011100" =>  data <= "00000000";  -- 51C = 0
      when "010100011101" =>  data <= "00000010";  -- 51D = 2
      when "010100011110" =>  data <= "01101001";  -- 51E = 69
      when "010100011111" =>  data <= "00000111";  -- 51F = 7
      when "010100100000" =>  data <= "11001000";  -- 520 = C8
      when "010100100001" =>  data <= "10011001";  -- 521 = 99
      when "010100100010" =>  data <= "00000000";  -- 522 = 0
      when "010100100011" =>  data <= "00000010";  -- 523 = 2
      when "010100100100" =>  data <= "01101001";  -- 524 = 69
      when "010100100101" =>  data <= "00000111";  -- 525 = 7
      when "010100100110" =>  data <= "11001000";  -- 526 = C8
      when "010100100111" =>  data <= "10011001";  -- 527 = 99
      when "010100101000" =>  data <= "00000000";  -- 528 = 0
      when "010100101001" =>  data <= "00000010";  -- 529 = 2
      when "010100101010" =>  data <= "10100000";  -- 52A = A0
      when "010100101011" =>  data <= "00000000";  -- 52B = 0
      when "010100101100" =>  data <= "00011000";  -- 52C = 18
      when "010100101101" =>  data <= "10111001";  -- 52D = B9
      when "010100101110" =>  data <= "00000000";  -- 52E = 0
      when "010100101111" =>  data <= "00000010";  -- 52F = 2
      when "010100110000" =>  data <= "11001001";  -- 530 = C9
      when "010100110001" =>  data <= "00000011";  -- 531 = 3
      when "010100110010" =>  data <= "11010000";  -- 532 = D0
      when "010100110011" =>  data <= "00110011";  -- 533 = 33
      when "010100110100" =>  data <= "11001000";  -- 534 = C8
      when "010100110101" =>  data <= "10111001";  -- 535 = B9
      when "010100110110" =>  data <= "00000000";  -- 536 = 0
      when "010100110111" =>  data <= "00000010";  -- 537 = 2
      when "010100111000" =>  data <= "11001001";  -- 538 = C9
      when "010100111001" =>  data <= "00001010";  -- 539 = A
      when "010100111010" =>  data <= "11010000";  -- 53A = D0
      when "010100111011" =>  data <= "00101011";  -- 53B = 2B
      when "010100111100" =>  data <= "11001000";  -- 53C = C8
      when "010100111101" =>  data <= "10111001";  -- 53D = B9
      when "010100111110" =>  data <= "00000000";  -- 53E = 0
      when "010100111111" =>  data <= "00000010";  -- 53F = 2
      when "010101000000" =>  data <= "11001001";  -- 540 = C9
      when "010101000001" =>  data <= "00010001";  -- 541 = 11
      when "010101000010" =>  data <= "11010000";  -- 542 = D0
      when "010101000011" =>  data <= "00100011";  -- 543 = 23
      when "010101000100" =>  data <= "11001000";  -- 544 = C8
      when "010101000101" =>  data <= "10111001";  -- 545 = B9
      when "010101000110" =>  data <= "00000000";  -- 546 = 0
      when "010101000111" =>  data <= "00000010";  -- 547 = 2
      when "010101001000" =>  data <= "11001001";  -- 548 = C9
      when "010101001001" =>  data <= "00011000";  -- 549 = 18
      when "010101001010" =>  data <= "11010000";  -- 54A = D0
      when "010101001011" =>  data <= "00011011";  -- 54B = 1B
      when "010101001100" =>  data <= "11001000";  -- 54C = C8
      when "010101001101" =>  data <= "10111001";  -- 54D = B9
      when "010101001110" =>  data <= "00000000";  -- 54E = 0
      when "010101001111" =>  data <= "00000010";  -- 54F = 2
      when "010101010000" =>  data <= "11001001";  -- 550 = C9
      when "010101010001" =>  data <= "00011111";  -- 551 = 1F
      when "010101010010" =>  data <= "11010000";  -- 552 = D0
      when "010101010011" =>  data <= "00010011";  -- 553 = 13
      when "010101010100" =>  data <= "11001000";  -- 554 = C8
      when "010101010101" =>  data <= "10111001";  -- 555 = B9
      when "010101010110" =>  data <= "00000000";  -- 556 = 0
      when "010101010111" =>  data <= "00000010";  -- 557 = 2
      when "010101011000" =>  data <= "11001001";  -- 558 = C9
      when "010101011001" =>  data <= "00100110";  -- 559 = 26
      when "010101011010" =>  data <= "11010000";  -- 55A = D0
      when "010101011011" =>  data <= "00001011";  -- 55B = B
      when "010101011100" =>  data <= "11001000";  -- 55C = C8
      when "010101011101" =>  data <= "10111001";  -- 55D = B9
      when "010101011110" =>  data <= "00000000";  -- 55E = 0
      when "010101011111" =>  data <= "00000010";  -- 55F = 2
      when "010101100000" =>  data <= "11001001";  -- 560 = C9
      when "010101100001" =>  data <= "00101101";  -- 561 = 2D
      when "010101100010" =>  data <= "11010000";  -- 562 = D0
      when "010101100011" =>  data <= "00000011";  -- 563 = 3
      when "010101100100" =>  data <= "01001100";  -- 564 = 4C
      when "010101100101" =>  data <= "01101100";  -- 565 = 6C
      when "010101100110" =>  data <= "11110101";  -- 566 = F5
      when "010101100111" =>  data <= "10101001";  -- 567 = A9
      when "010101101000" =>  data <= "01010000";  -- 568 = 50
      when "010101101001" =>  data <= "01001100";  -- 569 = 4C
      when "010101101010" =>  data <= "01000001";  -- 56A = 41
      when "010101101011" =>  data <= "11111001";  -- 56B = F9
      when "010101101100" =>  data <= "10101001";  -- 56C = A9
      when "010101101101" =>  data <= "00110100";  -- 56D = 34
      when "010101101110" =>  data <= "10001101";  -- 56E = 8D
      when "010101101111" =>  data <= "00000001";  -- 56F = 1
      when "010101110000" =>  data <= "10000000";  -- 570 = 80
      when "010101110001" =>  data <= "10101001";  -- 571 = A9
      when "010101110010" =>  data <= "01010010";  -- 572 = 52
      when "010101110011" =>  data <= "10001101";  -- 573 = 8D
      when "010101110100" =>  data <= "00000000";  -- 574 = 0
      when "010101110101" =>  data <= "00000010";  -- 575 = 2
      when "010101110110" =>  data <= "10101001";  -- 576 = A9
      when "010101110111" =>  data <= "00100100";  -- 577 = 24
      when "010101111000" =>  data <= "10001101";  -- 578 = 8D
      when "010101111001" =>  data <= "00000001";  -- 579 = 1
      when "010101111010" =>  data <= "00000010";  -- 57A = 2
      when "010101111011" =>  data <= "10101001";  -- 57B = A9
      when "010101111100" =>  data <= "01111000";  -- 57C = 78
      when "010101111101" =>  data <= "10001101";  -- 57D = 8D
      when "010101111110" =>  data <= "00000010";  -- 57E = 2
      when "010101111111" =>  data <= "00000010";  -- 57F = 2
      when "010110000000" =>  data <= "10101001";  -- 580 = A9
      when "010110000001" =>  data <= "00000000";  -- 581 = 0
      when "010110000010" =>  data <= "10100010";  -- 582 = A2
      when "010110000011" =>  data <= "00000000";  -- 583 = 0
      when "010110000100" =>  data <= "00011000";  -- 584 = 18
      when "010110000101" =>  data <= "01111101";  -- 585 = 7D
      when "010110000110" =>  data <= "00000000";  -- 586 = 0
      when "010110000111" =>  data <= "00000010";  -- 587 = 2
      when "010110001000" =>  data <= "00011000";  -- 588 = 18
      when "010110001001" =>  data <= "11101000";  -- 589 = E8
      when "010110001010" =>  data <= "01111101";  -- 58A = 7D
      when "010110001011" =>  data <= "00000000";  -- 58B = 0
      when "010110001100" =>  data <= "00000010";  -- 58C = 2
      when "010110001101" =>  data <= "00011000";  -- 58D = 18
      when "010110001110" =>  data <= "11101000";  -- 58E = E8
      when "010110001111" =>  data <= "01111101";  -- 58F = 7D
      when "010110010000" =>  data <= "00000000";  -- 590 = 0
      when "010110010001" =>  data <= "00000010";  -- 591 = 2
      when "010110010010" =>  data <= "11001001";  -- 592 = C9
      when "010110010011" =>  data <= "11101110";  -- 593 = EE
      when "010110010100" =>  data <= "11110000";  -- 594 = F0
      when "010110010101" =>  data <= "00000101";  -- 595 = 5
      when "010110010110" =>  data <= "10101001";  -- 596 = A9
      when "010110010111" =>  data <= "01010001";  -- 597 = 51
      when "010110011000" =>  data <= "01001100";  -- 598 = 4C
      when "010110011001" =>  data <= "01000001";  -- 599 = 41
      when "010110011010" =>  data <= "11111001";  -- 59A = F9
      when "010110011011" =>  data <= "10101001";  -- 59B = A9
      when "010110011100" =>  data <= "00110101";  -- 59C = 35
      when "010110011101" =>  data <= "10001101";  -- 59D = 8D
      when "010110011110" =>  data <= "00000001";  -- 59E = 1
      when "010110011111" =>  data <= "10000000";  -- 59F = 80
      when "010110100000" =>  data <= "10101001";  -- 5A0 = A9
      when "010110100001" =>  data <= "01101000";  -- 5A1 = 68
      when "010110100010" =>  data <= "10001101";  -- 5A2 = 8D
      when "010110100011" =>  data <= "00000000";  -- 5A3 = 0
      when "010110100100" =>  data <= "00000010";  -- 5A4 = 2
      when "010110100101" =>  data <= "10101001";  -- 5A5 = A9
      when "010110100110" =>  data <= "00010011";  -- 5A6 = 13
      when "010110100111" =>  data <= "10001101";  -- 5A7 = 8D
      when "010110101000" =>  data <= "00000001";  -- 5A8 = 1
      when "010110101001" =>  data <= "00000010";  -- 5A9 = 2
      when "010110101010" =>  data <= "10101001";  -- 5AA = A9
      when "010110101011" =>  data <= "10010101";  -- 5AB = 95
      when "010110101100" =>  data <= "10001101";  -- 5AC = 8D
      when "010110101101" =>  data <= "00000010";  -- 5AD = 2
      when "010110101110" =>  data <= "00000010";  -- 5AE = 2
      when "010110101111" =>  data <= "10101001";  -- 5AF = A9
      when "010110110000" =>  data <= "00000000";  -- 5B0 = 0
      when "010110110001" =>  data <= "10100000";  -- 5B1 = A0
      when "010110110010" =>  data <= "00000000";  -- 5B2 = 0
      when "010110110011" =>  data <= "00011000";  -- 5B3 = 18
      when "010110110100" =>  data <= "01111001";  -- 5B4 = 79
      when "010110110101" =>  data <= "00000000";  -- 5B5 = 0
      when "010110110110" =>  data <= "00000010";  -- 5B6 = 2
      when "010110110111" =>  data <= "00011000";  -- 5B7 = 18
      when "010110111000" =>  data <= "11001000";  -- 5B8 = C8
      when "010110111001" =>  data <= "01111001";  -- 5B9 = 79
      when "010110111010" =>  data <= "00000000";  -- 5BA = 0
      when "010110111011" =>  data <= "00000010";  -- 5BB = 2
      when "010110111100" =>  data <= "00011000";  -- 5BC = 18
      when "010110111101" =>  data <= "11001000";  -- 5BD = C8
      when "010110111110" =>  data <= "01111001";  -- 5BE = 79
      when "010110111111" =>  data <= "00000000";  -- 5BF = 0
      when "010111000000" =>  data <= "00000010";  -- 5C0 = 2
      when "010111000001" =>  data <= "11001001";  -- 5C1 = C9
      when "010111000010" =>  data <= "00010000";  -- 5C2 = 10
      when "010111000011" =>  data <= "11110000";  -- 5C3 = F0
      when "010111000100" =>  data <= "00000101";  -- 5C4 = 5
      when "010111000101" =>  data <= "10101001";  -- 5C5 = A9
      when "010111000110" =>  data <= "01010010";  -- 5C6 = 52
      when "010111000111" =>  data <= "01001100";  -- 5C7 = 4C
      when "010111001000" =>  data <= "01000001";  -- 5C8 = 41
      when "010111001001" =>  data <= "11111001";  -- 5C9 = F9
      when "010111001010" =>  data <= "10101001";  -- 5CA = A9
      when "010111001011" =>  data <= "00110110";  -- 5CB = 36
      when "010111001100" =>  data <= "10001101";  -- 5CC = 8D
      when "010111001101" =>  data <= "00000001";  -- 5CD = 1
      when "010111001110" =>  data <= "10000000";  -- 5CE = 80
      when "010111001111" =>  data <= "10101001";  -- 5CF = A9
      when "010111010000" =>  data <= "00110100";  -- 5D0 = 34
      when "010111010001" =>  data <= "10001101";  -- 5D1 = 8D
      when "010111010010" =>  data <= "00000000";  -- 5D2 = 0
      when "010111010011" =>  data <= "00000010";  -- 5D3 = 2
      when "010111010100" =>  data <= "10101001";  -- 5D4 = A9
      when "010111010101" =>  data <= "01010100";  -- 5D5 = 54
      when "010111010110" =>  data <= "10001101";  -- 5D6 = 8D
      when "010111010111" =>  data <= "00000001";  -- 5D7 = 1
      when "010111011000" =>  data <= "00000010";  -- 5D8 = 2
      when "010111011001" =>  data <= "10101001";  -- 5D9 = A9
      when "010111011010" =>  data <= "10010111";  -- 5DA = 97
      when "010111011011" =>  data <= "10001101";  -- 5DB = 8D
      when "010111011100" =>  data <= "00000010";  -- 5DC = 2
      when "010111011101" =>  data <= "00000010";  -- 5DD = 2
      when "010111011110" =>  data <= "10101001";  -- 5DE = A9
      when "010111011111" =>  data <= "11111111";  -- 5DF = FF
      when "010111100000" =>  data <= "10100000";  -- 5E0 = A0
      when "010111100001" =>  data <= "00000000";  -- 5E1 = 0
      when "010111100010" =>  data <= "00111001";  -- 5E2 = 39
      when "010111100011" =>  data <= "00000000";  -- 5E3 = 0
      when "010111100100" =>  data <= "00000010";  -- 5E4 = 2
      when "010111100101" =>  data <= "11001000";  -- 5E5 = C8
      when "010111100110" =>  data <= "00111001";  -- 5E6 = 39
      when "010111100111" =>  data <= "00000000";  -- 5E7 = 0
      when "010111101000" =>  data <= "00000010";  -- 5E8 = 2
      when "010111101001" =>  data <= "11001000";  -- 5E9 = C8
      when "010111101010" =>  data <= "00111001";  -- 5EA = 39
      when "010111101011" =>  data <= "00000000";  -- 5EB = 0
      when "010111101100" =>  data <= "00000010";  -- 5EC = 2
      when "010111101101" =>  data <= "11001001";  -- 5ED = C9
      when "010111101110" =>  data <= "00010100";  -- 5EE = 14
      when "010111101111" =>  data <= "11110000";  -- 5EF = F0
      when "010111110000" =>  data <= "00000101";  -- 5F0 = 5
      when "010111110001" =>  data <= "10101001";  -- 5F1 = A9
      when "010111110010" =>  data <= "01010011";  -- 5F2 = 53
      when "010111110011" =>  data <= "01001100";  -- 5F3 = 4C
      when "010111110100" =>  data <= "01000001";  -- 5F4 = 41
      when "010111110101" =>  data <= "11111001";  -- 5F5 = F9
      when "010111110110" =>  data <= "10101001";  -- 5F6 = A9
      when "010111110111" =>  data <= "00110111";  -- 5F7 = 37
      when "010111111000" =>  data <= "10001101";  -- 5F8 = 8D
      when "010111111001" =>  data <= "00000001";  -- 5F9 = 1
      when "010111111010" =>  data <= "10000000";  -- 5FA = 80
      when "010111111011" =>  data <= "10101001";  -- 5FB = A9
      when "010111111100" =>  data <= "00110100";  -- 5FC = 34
      when "010111111101" =>  data <= "10001101";  -- 5FD = 8D
      when "010111111110" =>  data <= "00000000";  -- 5FE = 0
      when "010111111111" =>  data <= "00000010";  -- 5FF = 2
      when "011000000000" =>  data <= "10101001";  -- 600 = A9
      when "011000000001" =>  data <= "01010100";  -- 601 = 54
      when "011000000010" =>  data <= "10001101";  -- 602 = 8D
      when "011000000011" =>  data <= "00000001";  -- 603 = 1
      when "011000000100" =>  data <= "00000010";  -- 604 = 2
      when "011000000101" =>  data <= "10101001";  -- 605 = A9
      when "011000000110" =>  data <= "10010111";  -- 606 = 97
      when "011000000111" =>  data <= "10001101";  -- 607 = 8D
      when "011000001000" =>  data <= "00000010";  -- 608 = 2
      when "011000001001" =>  data <= "00000010";  -- 609 = 2
      when "011000001010" =>  data <= "10101001";  -- 60A = A9
      when "011000001011" =>  data <= "11111111";  -- 60B = FF
      when "011000001100" =>  data <= "10100010";  -- 60C = A2
      when "011000001101" =>  data <= "00000000";  -- 60D = 0
      when "011000001110" =>  data <= "00111101";  -- 60E = 3D
      when "011000001111" =>  data <= "00000000";  -- 60F = 0
      when "011000010000" =>  data <= "00000010";  -- 610 = 2
      when "011000010001" =>  data <= "11101000";  -- 611 = E8
      when "011000010010" =>  data <= "00111101";  -- 612 = 3D
      when "011000010011" =>  data <= "00000000";  -- 613 = 0
      when "011000010100" =>  data <= "00000010";  -- 614 = 2
      when "011000010101" =>  data <= "11101000";  -- 615 = E8
      when "011000010110" =>  data <= "00111101";  -- 616 = 3D
      when "011000010111" =>  data <= "00000000";  -- 617 = 0
      when "011000011000" =>  data <= "00000010";  -- 618 = 2
      when "011000011001" =>  data <= "11001001";  -- 619 = C9
      when "011000011010" =>  data <= "00010100";  -- 61A = 14
      when "011000011011" =>  data <= "11110000";  -- 61B = F0
      when "011000011100" =>  data <= "00000101";  -- 61C = 5
      when "011000011101" =>  data <= "10101001";  -- 61D = A9
      when "011000011110" =>  data <= "01010100";  -- 61E = 54
      when "011000011111" =>  data <= "01001100";  -- 61F = 4C
      when "011000100000" =>  data <= "01000001";  -- 620 = 41
      when "011000100001" =>  data <= "11111001";  -- 621 = F9
      when "011000100010" =>  data <= "10101001";  -- 622 = A9
      when "011000100011" =>  data <= "00111000";  -- 623 = 38
      when "011000100100" =>  data <= "10001101";  -- 624 = 8D
      when "011000100101" =>  data <= "00000001";  -- 625 = 1
      when "011000100110" =>  data <= "10000000";  -- 626 = 80
      when "011000100111" =>  data <= "10101001";  -- 627 = A9
      when "011000101000" =>  data <= "01100100";  -- 628 = 64
      when "011000101001" =>  data <= "10000101";  -- 629 = 85
      when "011000101010" =>  data <= "00000000";  -- 62A = 0
      when "011000101011" =>  data <= "10101001";  -- 62B = A9
      when "011000101100" =>  data <= "00111001";  -- 62C = 39
      when "011000101101" =>  data <= "00011000";  -- 62D = 18
      when "011000101110" =>  data <= "01100101";  -- 62E = 65
      when "011000101111" =>  data <= "00000000";  -- 62F = 0
      when "011000110000" =>  data <= "11001001";  -- 630 = C9
      when "011000110001" =>  data <= "10011101";  -- 631 = 9D
      when "011000110010" =>  data <= "11110000";  -- 632 = F0
      when "011000110011" =>  data <= "00000101";  -- 633 = 5
      when "011000110100" =>  data <= "10101001";  -- 634 = A9
      when "011000110101" =>  data <= "01010101";  -- 635 = 55
      when "011000110110" =>  data <= "01001100";  -- 636 = 4C
      when "011000110111" =>  data <= "01000001";  -- 637 = 41
      when "011000111000" =>  data <= "11111001";  -- 638 = F9
      when "011000111001" =>  data <= "10101001";  -- 639 = A9
      when "011000111010" =>  data <= "00111001";  -- 63A = 39
      when "011000111011" =>  data <= "10001101";  -- 63B = 8D
      when "011000111100" =>  data <= "00000001";  -- 63C = 1
      when "011000111101" =>  data <= "10000000";  -- 63D = 80
      when "011000111110" =>  data <= "10101001";  -- 63E = A9
      when "011000111111" =>  data <= "10010101";  -- 63F = 95
      when "011001000000" =>  data <= "10000101";  -- 640 = 85
      when "011001000001" =>  data <= "00000000";  -- 641 = 0
      when "011001000010" =>  data <= "10101001";  -- 642 = A9
      when "011001000011" =>  data <= "01110110";  -- 643 = 76
      when "011001000100" =>  data <= "10000101";  -- 644 = 85
      when "011001000101" =>  data <= "00000001";  -- 645 = 1
      when "011001000110" =>  data <= "10101001";  -- 646 = A9
      when "011001000111" =>  data <= "01000101";  -- 647 = 45
      when "011001001000" =>  data <= "10000101";  -- 648 = 85
      when "011001001001" =>  data <= "00000010";  -- 649 = 2
      when "011001001010" =>  data <= "10100010";  -- 64A = A2
      when "011001001011" =>  data <= "00000000";  -- 64B = 0
      when "011001001100" =>  data <= "10101001";  -- 64C = A9
      when "011001001101" =>  data <= "00000000";  -- 64D = 0
      when "011001001110" =>  data <= "00011000";  -- 64E = 18
      when "011001001111" =>  data <= "01110101";  -- 64F = 75
      when "011001010000" =>  data <= "00000000";  -- 650 = 0
      when "011001010001" =>  data <= "11101000";  -- 651 = E8
      when "011001010010" =>  data <= "00011000";  -- 652 = 18
      when "011001010011" =>  data <= "01110101";  -- 653 = 75
      when "011001010100" =>  data <= "00000000";  -- 654 = 0
      when "011001010101" =>  data <= "11101000";  -- 655 = E8
      when "011001010110" =>  data <= "00011000";  -- 656 = 18
      when "011001010111" =>  data <= "01110101";  -- 657 = 75
      when "011001011000" =>  data <= "00000000";  -- 658 = 0
      when "011001011001" =>  data <= "11001001";  -- 659 = C9
      when "011001011010" =>  data <= "01010000";  -- 65A = 50
      when "011001011011" =>  data <= "11110000";  -- 65B = F0
      when "011001011100" =>  data <= "00000101";  -- 65C = 5
      when "011001011101" =>  data <= "10101001";  -- 65D = A9
      when "011001011110" =>  data <= "01010110";  -- 65E = 56
      when "011001011111" =>  data <= "01001100";  -- 65F = 4C
      when "011001100000" =>  data <= "01000001";  -- 660 = 41
      when "011001100001" =>  data <= "11111001";  -- 661 = F9
      when "011001100010" =>  data <= "10101001";  -- 662 = A9
      when "011001100011" =>  data <= "00111010";  -- 663 = 3A
      when "011001100100" =>  data <= "10001101";  -- 664 = 8D
      when "011001100101" =>  data <= "00000001";  -- 665 = 1
      when "011001100110" =>  data <= "10000000";  -- 666 = 80
      when "011001100111" =>  data <= "10101001";  -- 667 = A9
      when "011001101000" =>  data <= "01100100";  -- 668 = 64
      when "011001101001" =>  data <= "10000101";  -- 669 = 85
      when "011001101010" =>  data <= "00000000";  -- 66A = 0
      when "011001101011" =>  data <= "10101001";  -- 66B = A9
      when "011001101100" =>  data <= "00111001";  -- 66C = 39
      when "011001101101" =>  data <= "00100101";  -- 66D = 25
      when "011001101110" =>  data <= "00000000";  -- 66E = 0
      when "011001101111" =>  data <= "11001001";  -- 66F = C9
      when "011001110000" =>  data <= "00100000";  -- 670 = 20
      when "011001110001" =>  data <= "11110000";  -- 671 = F0
      when "011001110010" =>  data <= "00000101";  -- 672 = 5
      when "011001110011" =>  data <= "10101001";  -- 673 = A9
      when "011001110100" =>  data <= "01010111";  -- 674 = 57
      when "011001110101" =>  data <= "01001100";  -- 675 = 4C
      when "011001110110" =>  data <= "01000001";  -- 676 = 41
      when "011001110111" =>  data <= "11111001";  -- 677 = F9
      when "011001111000" =>  data <= "10101001";  -- 678 = A9
      when "011001111001" =>  data <= "00111011";  -- 679 = 3B
      when "011001111010" =>  data <= "10001101";  -- 67A = 8D
      when "011001111011" =>  data <= "00000001";  -- 67B = 1
      when "011001111100" =>  data <= "10000000";  -- 67C = 80
      when "011001111101" =>  data <= "10101001";  -- 67D = A9
      when "011001111110" =>  data <= "10010101";  -- 67E = 95
      when "011001111111" =>  data <= "10000101";  -- 67F = 85
      when "011010000000" =>  data <= "00000000";  -- 680 = 0
      when "011010000001" =>  data <= "10101001";  -- 681 = A9
      when "011010000010" =>  data <= "01110110";  -- 682 = 76
      when "011010000011" =>  data <= "10000101";  -- 683 = 85
      when "011010000100" =>  data <= "00000001";  -- 684 = 1
      when "011010000101" =>  data <= "10101001";  -- 685 = A9
      when "011010000110" =>  data <= "01000101";  -- 686 = 45
      when "011010000111" =>  data <= "10000101";  -- 687 = 85
      when "011010001000" =>  data <= "00000010";  -- 688 = 2
      when "011010001001" =>  data <= "10100010";  -- 689 = A2
      when "011010001010" =>  data <= "00000000";  -- 68A = 0
      when "011010001011" =>  data <= "10101001";  -- 68B = A9
      when "011010001100" =>  data <= "11111111";  -- 68C = FF
      when "011010001101" =>  data <= "00110101";  -- 68D = 35
      when "011010001110" =>  data <= "00000000";  -- 68E = 0
      when "011010001111" =>  data <= "11101000";  -- 68F = E8
      when "011010010000" =>  data <= "00110101";  -- 690 = 35
      when "011010010001" =>  data <= "00000000";  -- 691 = 0
      when "011010010010" =>  data <= "11101000";  -- 692 = E8
      when "011010010011" =>  data <= "00110101";  -- 693 = 35
      when "011010010100" =>  data <= "00000000";  -- 694 = 0
      when "011010010101" =>  data <= "11001001";  -- 695 = C9
      when "011010010110" =>  data <= "00000100";  -- 696 = 4
      when "011010010111" =>  data <= "11110000";  -- 697 = F0
      when "011010011000" =>  data <= "00000101";  -- 698 = 5
      when "011010011001" =>  data <= "10101001";  -- 699 = A9
      when "011010011010" =>  data <= "01011000";  -- 69A = 58
      when "011010011011" =>  data <= "01001100";  -- 69B = 4C
      when "011010011100" =>  data <= "01000001";  -- 69C = 41
      when "011010011101" =>  data <= "11111001";  -- 69D = F9
      when "011010011110" =>  data <= "10101001";  -- 69E = A9
      when "011010011111" =>  data <= "00111100";  -- 69F = 3C
      when "011010100000" =>  data <= "10001101";  -- 6A0 = 8D
      when "011010100001" =>  data <= "00000001";  -- 6A1 = 1
      when "011010100010" =>  data <= "10000000";  -- 6A2 = 80
      when "011010100011" =>  data <= "10101001";  -- 6A3 = A9
      when "011010100100" =>  data <= "10010111";  -- 6A4 = 97
      when "011010100101" =>  data <= "10001101";  -- 6A5 = 8D
      when "011010100110" =>  data <= "00000000";  -- 6A6 = 0
      when "011010100111" =>  data <= "00000010";  -- 6A7 = 2
      when "011010101000" =>  data <= "10101001";  -- 6A8 = A9
      when "011010101001" =>  data <= "01111000";  -- 6A9 = 78
      when "011010101010" =>  data <= "10001101";  -- 6AA = 8D
      when "011010101011" =>  data <= "00000001";  -- 6AB = 1
      when "011010101100" =>  data <= "00000010";  -- 6AC = 2
      when "011010101101" =>  data <= "10101001";  -- 6AD = A9
      when "011010101110" =>  data <= "01000101";  -- 6AE = 45
      when "011010101111" =>  data <= "10001101";  -- 6AF = 8D
      when "011010110000" =>  data <= "00000010";  -- 6B0 = 2
      when "011010110001" =>  data <= "00000010";  -- 6B1 = 2
      when "011010110010" =>  data <= "10100010";  -- 6B2 = A2
      when "011010110011" =>  data <= "00000000";  -- 6B3 = 0
      when "011010110100" =>  data <= "10101001";  -- 6B4 = A9
      when "011010110101" =>  data <= "10010111";  -- 6B5 = 97
      when "011010110110" =>  data <= "11011101";  -- 6B6 = DD
      when "011010110111" =>  data <= "00000000";  -- 6B7 = 0
      when "011010111000" =>  data <= "00000010";  -- 6B8 = 2
      when "011010111001" =>  data <= "11010000";  -- 6B9 = D0
      when "011010111010" =>  data <= "00010011";  -- 6BA = 13
      when "011010111011" =>  data <= "10101001";  -- 6BB = A9
      when "011010111100" =>  data <= "01111000";  -- 6BC = 78
      when "011010111101" =>  data <= "11101000";  -- 6BD = E8
      when "011010111110" =>  data <= "11011101";  -- 6BE = DD
      when "011010111111" =>  data <= "00000000";  -- 6BF = 0
      when "011011000000" =>  data <= "00000010";  -- 6C0 = 2
      when "011011000001" =>  data <= "11010000";  -- 6C1 = D0
      when "011011000010" =>  data <= "00001011";  -- 6C2 = B
      when "011011000011" =>  data <= "10101001";  -- 6C3 = A9
      when "011011000100" =>  data <= "01000101";  -- 6C4 = 45
      when "011011000101" =>  data <= "11101000";  -- 6C5 = E8
      when "011011000110" =>  data <= "11011101";  -- 6C6 = DD
      when "011011000111" =>  data <= "00000000";  -- 6C7 = 0
      when "011011001000" =>  data <= "00000010";  -- 6C8 = 2
      when "011011001001" =>  data <= "11010000";  -- 6C9 = D0
      when "011011001010" =>  data <= "00000011";  -- 6CA = 3
      when "011011001011" =>  data <= "01001100";  -- 6CB = 4C
      when "011011001100" =>  data <= "11010011";  -- 6CC = D3
      when "011011001101" =>  data <= "11110110";  -- 6CD = F6
      when "011011001110" =>  data <= "10101001";  -- 6CE = A9
      when "011011001111" =>  data <= "01011001";  -- 6CF = 59
      when "011011010000" =>  data <= "01001100";  -- 6D0 = 4C
      when "011011010001" =>  data <= "01000001";  -- 6D1 = 41
      when "011011010010" =>  data <= "11111001";  -- 6D2 = F9
      when "011011010011" =>  data <= "10101001";  -- 6D3 = A9
      when "011011010100" =>  data <= "00111101";  -- 6D4 = 3D
      when "011011010101" =>  data <= "10001101";  -- 6D5 = 8D
      when "011011010110" =>  data <= "00000001";  -- 6D6 = 1
      when "011011010111" =>  data <= "10000000";  -- 6D7 = 80
      when "011011011000" =>  data <= "10101001";  -- 6D8 = A9
      when "011011011001" =>  data <= "10010111";  -- 6D9 = 97
      when "011011011010" =>  data <= "10001101";  -- 6DA = 8D
      when "011011011011" =>  data <= "00000000";  -- 6DB = 0
      when "011011011100" =>  data <= "00000010";  -- 6DC = 2
      when "011011011101" =>  data <= "10101001";  -- 6DD = A9
      when "011011011110" =>  data <= "01111000";  -- 6DE = 78
      when "011011011111" =>  data <= "10001101";  -- 6DF = 8D
      when "011011100000" =>  data <= "00000001";  -- 6E0 = 1
      when "011011100001" =>  data <= "00000010";  -- 6E1 = 2
      when "011011100010" =>  data <= "10101001";  -- 6E2 = A9
      when "011011100011" =>  data <= "01000101";  -- 6E3 = 45
      when "011011100100" =>  data <= "10001101";  -- 6E4 = 8D
      when "011011100101" =>  data <= "00000010";  -- 6E5 = 2
      when "011011100110" =>  data <= "00000010";  -- 6E6 = 2
      when "011011100111" =>  data <= "10100000";  -- 6E7 = A0
      when "011011101000" =>  data <= "00000000";  -- 6E8 = 0
      when "011011101001" =>  data <= "10101001";  -- 6E9 = A9
      when "011011101010" =>  data <= "10010111";  -- 6EA = 97
      when "011011101011" =>  data <= "11011001";  -- 6EB = D9
      when "011011101100" =>  data <= "00000000";  -- 6EC = 0
      when "011011101101" =>  data <= "00000010";  -- 6ED = 2
      when "011011101110" =>  data <= "11010000";  -- 6EE = D0
      when "011011101111" =>  data <= "00010011";  -- 6EF = 13
      when "011011110000" =>  data <= "10101001";  -- 6F0 = A9
      when "011011110001" =>  data <= "01111000";  -- 6F1 = 78
      when "011011110010" =>  data <= "11001000";  -- 6F2 = C8
      when "011011110011" =>  data <= "11011001";  -- 6F3 = D9
      when "011011110100" =>  data <= "00000000";  -- 6F4 = 0
      when "011011110101" =>  data <= "00000010";  -- 6F5 = 2
      when "011011110110" =>  data <= "11010000";  -- 6F6 = D0
      when "011011110111" =>  data <= "00001011";  -- 6F7 = B
      when "011011111000" =>  data <= "10101001";  -- 6F8 = A9
      when "011011111001" =>  data <= "01000101";  -- 6F9 = 45
      when "011011111010" =>  data <= "11001000";  -- 6FA = C8
      when "011011111011" =>  data <= "11011001";  -- 6FB = D9
      when "011011111100" =>  data <= "00000000";  -- 6FC = 0
      when "011011111101" =>  data <= "00000010";  -- 6FD = 2
      when "011011111110" =>  data <= "11010000";  -- 6FE = D0
      when "011011111111" =>  data <= "00000011";  -- 6FF = 3
      when "011100000000" =>  data <= "01001100";  -- 700 = 4C
      when "011100000001" =>  data <= "00001000";  -- 701 = 8
      when "011100000010" =>  data <= "11110111";  -- 702 = F7
      when "011100000011" =>  data <= "10101001";  -- 703 = A9
      when "011100000100" =>  data <= "01011010";  -- 704 = 5A
      when "011100000101" =>  data <= "01001100";  -- 705 = 4C
      when "011100000110" =>  data <= "01000001";  -- 706 = 41
      when "011100000111" =>  data <= "11111001";  -- 707 = F9
      when "011100001000" =>  data <= "10101001";  -- 708 = A9
      when "011100001001" =>  data <= "00111110";  -- 709 = 3E
      when "011100001010" =>  data <= "10001101";  -- 70A = 8D
      when "011100001011" =>  data <= "00000001";  -- 70B = 1
      when "011100001100" =>  data <= "10000000";  -- 70C = 80
      when "011100001101" =>  data <= "10101001";  -- 70D = A9
      when "011100001110" =>  data <= "10010111";  -- 70E = 97
      when "011100001111" =>  data <= "10001101";  -- 70F = 8D
      when "011100010000" =>  data <= "00000000";  -- 710 = 0
      when "011100010001" =>  data <= "00000010";  -- 711 = 2
      when "011100010010" =>  data <= "10101001";  -- 712 = A9
      when "011100010011" =>  data <= "01111000";  -- 713 = 78
      when "011100010100" =>  data <= "10001101";  -- 714 = 8D
      when "011100010101" =>  data <= "00000001";  -- 715 = 1
      when "011100010110" =>  data <= "00000010";  -- 716 = 2
      when "011100010111" =>  data <= "10101001";  -- 717 = A9
      when "011100011000" =>  data <= "01000101";  -- 718 = 45
      when "011100011001" =>  data <= "10001101";  -- 719 = 8D
      when "011100011010" =>  data <= "00000010";  -- 71A = 2
      when "011100011011" =>  data <= "00000010";  -- 71B = 2
      when "011100011100" =>  data <= "10100010";  -- 71C = A2
      when "011100011101" =>  data <= "00000000";  -- 71D = 0
      when "011100011110" =>  data <= "10101001";  -- 71E = A9
      when "011100011111" =>  data <= "10010111";  -- 71F = 97
      when "011100100000" =>  data <= "11011101";  -- 720 = DD
      when "011100100001" =>  data <= "00000000";  -- 721 = 0
      when "011100100010" =>  data <= "00000010";  -- 722 = 2
      when "011100100011" =>  data <= "11010000";  -- 723 = D0
      when "011100100100" =>  data <= "00010011";  -- 724 = 13
      when "011100100101" =>  data <= "10101001";  -- 725 = A9
      when "011100100110" =>  data <= "01111000";  -- 726 = 78
      when "011100100111" =>  data <= "11101000";  -- 727 = E8
      when "011100101000" =>  data <= "11011101";  -- 728 = DD
      when "011100101001" =>  data <= "00000000";  -- 729 = 0
      when "011100101010" =>  data <= "00000010";  -- 72A = 2
      when "011100101011" =>  data <= "11010000";  -- 72B = D0
      when "011100101100" =>  data <= "00001011";  -- 72C = B
      when "011100101101" =>  data <= "10101001";  -- 72D = A9
      when "011100101110" =>  data <= "01000101";  -- 72E = 45
      when "011100101111" =>  data <= "11101000";  -- 72F = E8
      when "011100110000" =>  data <= "11011101";  -- 730 = DD
      when "011100110001" =>  data <= "00000000";  -- 731 = 0
      when "011100110010" =>  data <= "00000010";  -- 732 = 2
      when "011100110011" =>  data <= "11010000";  -- 733 = D0
      when "011100110100" =>  data <= "00000011";  -- 734 = 3
      when "011100110101" =>  data <= "01001100";  -- 735 = 4C
      when "011100110110" =>  data <= "00111101";  -- 736 = 3D
      when "011100110111" =>  data <= "11110111";  -- 737 = F7
      when "011100111000" =>  data <= "10101001";  -- 738 = A9
      when "011100111001" =>  data <= "01011011";  -- 739 = 5B
      when "011100111010" =>  data <= "01001100";  -- 73A = 4C
      when "011100111011" =>  data <= "01000001";  -- 73B = 41
      when "011100111100" =>  data <= "11111001";  -- 73C = F9
      when "011100111101" =>  data <= "10101001";  -- 73D = A9
      when "011100111110" =>  data <= "00111111";  -- 73E = 3F
      when "011100111111" =>  data <= "10001101";  -- 73F = 8D
      when "011101000000" =>  data <= "00000001";  -- 740 = 1
      when "011101000001" =>  data <= "10000000";  -- 741 = 80
      when "011101000010" =>  data <= "10101001";  -- 742 = A9
      when "011101000011" =>  data <= "10010101";  -- 743 = 95
      when "011101000100" =>  data <= "10000101";  -- 744 = 85
      when "011101000101" =>  data <= "00000010";  -- 745 = 2
      when "011101000110" =>  data <= "10101001";  -- 746 = A9
      when "011101000111" =>  data <= "00000000";  -- 747 = 0
      when "011101001000" =>  data <= "10101001";  -- 748 = A9
      when "011101001001" =>  data <= "10010101";  -- 749 = 95
      when "011101001010" =>  data <= "11000101";  -- 74A = C5
      when "011101001011" =>  data <= "00000010";  -- 74B = 2
      when "011101001100" =>  data <= "11110000";  -- 74C = F0
      when "011101001101" =>  data <= "00000101";  -- 74D = 5
      when "011101001110" =>  data <= "10101001";  -- 74E = A9
      when "011101001111" =>  data <= "01011100";  -- 74F = 5C
      when "011101010000" =>  data <= "01001100";  -- 750 = 4C
      when "011101010001" =>  data <= "01000001";  -- 751 = 41
      when "011101010010" =>  data <= "11111001";  -- 752 = F9
      when "011101010011" =>  data <= "10101001";  -- 753 = A9
      when "011101010100" =>  data <= "01110101";  -- 754 = 75
      when "011101010101" =>  data <= "10000101";  -- 755 = 85
      when "011101010110" =>  data <= "00000010";  -- 756 = 2
      when "011101010111" =>  data <= "10101001";  -- 757 = A9
      when "011101011000" =>  data <= "01100111";  -- 758 = 67
      when "011101011001" =>  data <= "11000101";  -- 759 = C5
      when "011101011010" =>  data <= "00000010";  -- 75A = 2
      when "011101011011" =>  data <= "11010000";  -- 75B = D0
      when "011101011100" =>  data <= "00000101";  -- 75C = 5
      when "011101011101" =>  data <= "10101001";  -- 75D = A9
      when "011101011110" =>  data <= "01011101";  -- 75E = 5D
      when "011101011111" =>  data <= "01001100";  -- 75F = 4C
      when "011101100000" =>  data <= "01000001";  -- 760 = 41
      when "011101100001" =>  data <= "11111001";  -- 761 = F9
      when "011101100010" =>  data <= "10101001";  -- 762 = A9
      when "011101100011" =>  data <= "01000000";  -- 763 = 40
      when "011101100100" =>  data <= "10001101";  -- 764 = 8D
      when "011101100101" =>  data <= "00000001";  -- 765 = 1
      when "011101100110" =>  data <= "10000000";  -- 766 = 80
      when "011101100111" =>  data <= "10101001";  -- 767 = A9
      when "011101101000" =>  data <= "00110110";  -- 768 = 36
      when "011101101001" =>  data <= "10000101";  -- 769 = 85
      when "011101101010" =>  data <= "00000010";  -- 76A = 2
      when "011101101011" =>  data <= "10101001";  -- 76B = A9
      when "011101101100" =>  data <= "00000000";  -- 76C = 0
      when "011101101101" =>  data <= "10100010";  -- 76D = A2
      when "011101101110" =>  data <= "00110110";  -- 76E = 36
      when "011101101111" =>  data <= "11100100";  -- 76F = E4
      when "011101110000" =>  data <= "00000010";  -- 770 = 2
      when "011101110001" =>  data <= "11110000";  -- 771 = F0
      when "011101110010" =>  data <= "00000101";  -- 772 = 5
      when "011101110011" =>  data <= "10101001";  -- 773 = A9
      when "011101110100" =>  data <= "01011110";  -- 774 = 5E
      when "011101110101" =>  data <= "01001100";  -- 775 = 4C
      when "011101110110" =>  data <= "01000001";  -- 776 = 41
      when "011101110111" =>  data <= "11111001";  -- 777 = F9
      when "011101111000" =>  data <= "10101001";  -- 778 = A9
      when "011101111001" =>  data <= "01010111";  -- 779 = 57
      when "011101111010" =>  data <= "10000101";  -- 77A = 85
      when "011101111011" =>  data <= "00000010";  -- 77B = 2
      when "011101111100" =>  data <= "10100010";  -- 77C = A2
      when "011101111101" =>  data <= "00111001";  -- 77D = 39
      when "011101111110" =>  data <= "11100100";  -- 77E = E4
      when "011101111111" =>  data <= "00000010";  -- 77F = 2
      when "011110000000" =>  data <= "11010000";  -- 780 = D0
      when "011110000001" =>  data <= "00000101";  -- 781 = 5
      when "011110000010" =>  data <= "10101001";  -- 782 = A9
      when "011110000011" =>  data <= "01011111";  -- 783 = 5F
      when "011110000100" =>  data <= "01001100";  -- 784 = 4C
      when "011110000101" =>  data <= "01000001";  -- 785 = 41
      when "011110000110" =>  data <= "11111001";  -- 786 = F9
      when "011110000111" =>  data <= "10101001";  -- 787 = A9
      when "011110001000" =>  data <= "01000001";  -- 788 = 41
      when "011110001001" =>  data <= "10001101";  -- 789 = 8D
      when "011110001010" =>  data <= "00000001";  -- 78A = 1
      when "011110001011" =>  data <= "10000000";  -- 78B = 80
      when "011110001100" =>  data <= "10101001";  -- 78C = A9
      when "011110001101" =>  data <= "01110101";  -- 78D = 75
      when "011110001110" =>  data <= "10000101";  -- 78E = 85
      when "011110001111" =>  data <= "00000010";  -- 78F = 2
      when "011110010000" =>  data <= "10101001";  -- 790 = A9
      when "011110010001" =>  data <= "00000000";  -- 791 = 0
      when "011110010010" =>  data <= "10100000";  -- 792 = A0
      when "011110010011" =>  data <= "01110101";  -- 793 = 75
      when "011110010100" =>  data <= "11000100";  -- 794 = C4
      when "011110010101" =>  data <= "00000010";  -- 795 = 2
      when "011110010110" =>  data <= "11110000";  -- 796 = F0
      when "011110010111" =>  data <= "00000101";  -- 797 = 5
      when "011110011000" =>  data <= "10101001";  -- 798 = A9
      when "011110011001" =>  data <= "01100000";  -- 799 = 60
      when "011110011010" =>  data <= "01001100";  -- 79A = 4C
      when "011110011011" =>  data <= "01000001";  -- 79B = 41
      when "011110011100" =>  data <= "11111001";  -- 79C = F9
      when "011110011101" =>  data <= "10101001";  -- 79D = A9
      when "011110011110" =>  data <= "01000011";  -- 79E = 43
      when "011110011111" =>  data <= "10000101";  -- 79F = 85
      when "011110100000" =>  data <= "00000010";  -- 7A0 = 2
      when "011110100001" =>  data <= "10100000";  -- 7A1 = A0
      when "011110100010" =>  data <= "00100100";  -- 7A2 = 24
      when "011110100011" =>  data <= "11000100";  -- 7A3 = C4
      when "011110100100" =>  data <= "00000010";  -- 7A4 = 2
      when "011110100101" =>  data <= "11010000";  -- 7A5 = D0
      when "011110100110" =>  data <= "00000101";  -- 7A6 = 5
      when "011110100111" =>  data <= "10101001";  -- 7A7 = A9
      when "011110101000" =>  data <= "01100001";  -- 7A8 = 61
      when "011110101001" =>  data <= "01001100";  -- 7A9 = 4C
      when "011110101010" =>  data <= "01000001";  -- 7AA = 41
      when "011110101011" =>  data <= "11111001";  -- 7AB = F9
      when "011110101100" =>  data <= "10101001";  -- 7AC = A9
      when "011110101101" =>  data <= "01000010";  -- 7AD = 42
      when "011110101110" =>  data <= "10001101";  -- 7AE = 8D
      when "011110101111" =>  data <= "00000001";  -- 7AF = 1
      when "011110110000" =>  data <= "10000000";  -- 7B0 = 80
      when "011110110001" =>  data <= "01011000";  -- 7B1 = 58
      when "011110110010" =>  data <= "10101001";  -- 7B2 = A9
      when "011110110011" =>  data <= "00000000";  -- 7B3 = 0
      when "011110110100" =>  data <= "10000101";  -- 7B4 = 85
      when "011110110101" =>  data <= "00000101";  -- 7B5 = 5
      when "011110110110" =>  data <= "10101001";  -- 7B6 = A9
      when "011110110111" =>  data <= "00000001";  -- 7B7 = 1
      when "011110111000" =>  data <= "10000101";  -- 7B8 = 85
      when "011110111001" =>  data <= "00000100";  -- 7B9 = 4
      when "011110111010" =>  data <= "10101001";  -- 7BA = A9
      when "011110111011" =>  data <= "00010000";  -- 7BB = 10
      when "011110111100" =>  data <= "10001101";  -- 7BC = 8D
      when "011110111101" =>  data <= "00000101";  -- 7BD = 5
      when "011110111110" =>  data <= "10000000";  -- 7BE = 80
      when "011110111111" =>  data <= "10001101";  -- 7BF = 8D
      when "011111000000" =>  data <= "00000100";  -- 7C0 = 4
      when "011111000001" =>  data <= "10000000";  -- 7C1 = 80
      when "011111000010" =>  data <= "10100010";  -- 7C2 = A2
      when "011111000011" =>  data <= "00000000";  -- 7C3 = 0
      when "011111000100" =>  data <= "11101000";  -- 7C4 = E8
      when "011111000101" =>  data <= "11101000";  -- 7C5 = E8
      when "011111000110" =>  data <= "11101000";  -- 7C6 = E8
      when "011111000111" =>  data <= "11101000";  -- 7C7 = E8
      when "011111001000" =>  data <= "11101000";  -- 7C8 = E8
      when "011111001001" =>  data <= "11101000";  -- 7C9 = E8
      when "011111001010" =>  data <= "11101000";  -- 7CA = E8
      when "011111001011" =>  data <= "11101000";  -- 7CB = E8
      when "011111001100" =>  data <= "11101000";  -- 7CC = E8
      when "011111001101" =>  data <= "11101000";  -- 7CD = E8
      when "011111001110" =>  data <= "11101000";  -- 7CE = E8
      when "011111001111" =>  data <= "11101000";  -- 7CF = E8
      when "011111010000" =>  data <= "11101000";  -- 7D0 = E8
      when "011111010001" =>  data <= "11101000";  -- 7D1 = E8
      when "011111010010" =>  data <= "11101000";  -- 7D2 = E8
      when "011111010011" =>  data <= "11101000";  -- 7D3 = E8
      when "011111010100" =>  data <= "11100000";  -- 7D4 = E0
      when "011111010101" =>  data <= "00010000";  -- 7D5 = 10
      when "011111010110" =>  data <= "11110000";  -- 7D6 = F0
      when "011111010111" =>  data <= "00000101";  -- 7D7 = 5
      when "011111011000" =>  data <= "10101001";  -- 7D8 = A9
      when "011111011001" =>  data <= "01100010";  -- 7D9 = 62
      when "011111011010" =>  data <= "01001100";  -- 7DA = 4C
      when "011111011011" =>  data <= "01000001";  -- 7DB = 41
      when "011111011100" =>  data <= "11111001";  -- 7DC = F9
      when "011111011101" =>  data <= "10100101";  -- 7DD = A5
      when "011111011110" =>  data <= "00000101";  -- 7DE = 5
      when "011111011111" =>  data <= "11001001";  -- 7DF = C9
      when "011111100000" =>  data <= "00000001";  -- 7E0 = 1
      when "011111100001" =>  data <= "11110000";  -- 7E1 = F0
      when "011111100010" =>  data <= "00000101";  -- 7E2 = 5
      when "011111100011" =>  data <= "10101001";  -- 7E3 = A9
      when "011111100100" =>  data <= "01100011";  -- 7E4 = 63
      when "011111100101" =>  data <= "01001100";  -- 7E5 = 4C
      when "011111100110" =>  data <= "01000001";  -- 7E6 = 41
      when "011111100111" =>  data <= "11111001";  -- 7E7 = F9
      when "011111101000" =>  data <= "01111000";  -- 7E8 = 78
      when "011111101001" =>  data <= "10101001";  -- 7E9 = A9
      when "011111101010" =>  data <= "00000000";  -- 7EA = 0
      when "011111101011" =>  data <= "10000101";  -- 7EB = 85
      when "011111101100" =>  data <= "00000101";  -- 7EC = 5
      when "011111101101" =>  data <= "10101001";  -- 7ED = A9
      when "011111101110" =>  data <= "00000001";  -- 7EE = 1
      when "011111101111" =>  data <= "10000101";  -- 7EF = 85
      when "011111110000" =>  data <= "00000100";  -- 7F0 = 4
      when "011111110001" =>  data <= "10101001";  -- 7F1 = A9
      when "011111110010" =>  data <= "00010000";  -- 7F2 = 10
      when "011111110011" =>  data <= "10001101";  -- 7F3 = 8D
      when "011111110100" =>  data <= "00000101";  -- 7F4 = 5
      when "011111110101" =>  data <= "10000000";  -- 7F5 = 80
      when "011111110110" =>  data <= "10001101";  -- 7F6 = 8D
      when "011111110111" =>  data <= "00000100";  -- 7F7 = 4
      when "011111111000" =>  data <= "10000000";  -- 7F8 = 80
      when "011111111001" =>  data <= "10100010";  -- 7F9 = A2
      when "011111111010" =>  data <= "00000000";  -- 7FA = 0
      when "011111111011" =>  data <= "11101000";  -- 7FB = E8
      when "011111111100" =>  data <= "11101000";  -- 7FC = E8
      when "011111111101" =>  data <= "11101000";  -- 7FD = E8
      when "011111111110" =>  data <= "11101000";  -- 7FE = E8
      when "011111111111" =>  data <= "11101000";  -- 7FF = E8
      when "100000000000" =>  data <= "11101000";  -- 800 = E8
      when "100000000001" =>  data <= "11101000";  -- 801 = E8
      when "100000000010" =>  data <= "11101000";  -- 802 = E8
      when "100000000011" =>  data <= "11101000";  -- 803 = E8
      when "100000000100" =>  data <= "11101000";  -- 804 = E8
      when "100000000101" =>  data <= "11101000";  -- 805 = E8
      when "100000000110" =>  data <= "11101000";  -- 806 = E8
      when "100000000111" =>  data <= "11101000";  -- 807 = E8
      when "100000001000" =>  data <= "11101000";  -- 808 = E8
      when "100000001001" =>  data <= "11101000";  -- 809 = E8
      when "100000001010" =>  data <= "11101000";  -- 80A = E8
      when "100000001011" =>  data <= "11100000";  -- 80B = E0
      when "100000001100" =>  data <= "00010000";  -- 80C = 10
      when "100000001101" =>  data <= "11110000";  -- 80D = F0
      when "100000001110" =>  data <= "00000101";  -- 80E = 5
      when "100000001111" =>  data <= "10101001";  -- 80F = A9
      when "100000010000" =>  data <= "01100010";  -- 810 = 62
      when "100000010001" =>  data <= "01001100";  -- 811 = 4C
      when "100000010010" =>  data <= "01000001";  -- 812 = 41
      when "100000010011" =>  data <= "11111001";  -- 813 = F9
      when "100000010100" =>  data <= "10100101";  -- 814 = A5
      when "100000010101" =>  data <= "00000101";  -- 815 = 5
      when "100000010110" =>  data <= "11001001";  -- 816 = C9
      when "100000010111" =>  data <= "00000000";  -- 817 = 0
      when "100000011000" =>  data <= "11110000";  -- 818 = F0
      when "100000011001" =>  data <= "00000101";  -- 819 = 5
      when "100000011010" =>  data <= "10101001";  -- 81A = A9
      when "100000011011" =>  data <= "01100011";  -- 81B = 63
      when "100000011100" =>  data <= "01001100";  -- 81C = 4C
      when "100000011101" =>  data <= "01000001";  -- 81D = 41
      when "100000011110" =>  data <= "11111001";  -- 81E = F9
      when "100000011111" =>  data <= "10101001";  -- 81F = A9
      when "100000100000" =>  data <= "00000000";  -- 820 = 0
      when "100000100001" =>  data <= "10000101";  -- 821 = 85
      when "100000100010" =>  data <= "00000100";  -- 822 = 4
      when "100000100011" =>  data <= "10001101";  -- 823 = 8D
      when "100000100100" =>  data <= "00000101";  -- 824 = 5
      when "100000100101" =>  data <= "10000000";  -- 825 = 80
      when "100000100110" =>  data <= "10101001";  -- 826 = A9
      when "100000100111" =>  data <= "01000011";  -- 827 = 43
      when "100000101000" =>  data <= "10001101";  -- 828 = 8D
      when "100000101001" =>  data <= "00000001";  -- 829 = 1
      when "100000101010" =>  data <= "10000000";  -- 82A = 80
      when "100000101011" =>  data <= "10101001";  -- 82B = A9
      when "100000101100" =>  data <= "00000000";  -- 82C = 0
      when "100000101101" =>  data <= "10000101";  -- 82D = 85
      when "100000101110" =>  data <= "00000111";  -- 82E = 7
      when "100000101111" =>  data <= "10101001";  -- 82F = A9
      when "100000110000" =>  data <= "00000001";  -- 830 = 1
      when "100000110001" =>  data <= "10000101";  -- 831 = 85
      when "100000110010" =>  data <= "00000110";  -- 832 = 6
      when "100000110011" =>  data <= "10101001";  -- 833 = A9
      when "100000110100" =>  data <= "00010000";  -- 834 = 10
      when "100000110101" =>  data <= "10001101";  -- 835 = 8D
      when "100000110110" =>  data <= "00000111";  -- 836 = 7
      when "100000110111" =>  data <= "10000000";  -- 837 = 80
      when "100000111000" =>  data <= "10001101";  -- 838 = 8D
      when "100000111001" =>  data <= "00000110";  -- 839 = 6
      when "100000111010" =>  data <= "10000000";  -- 83A = 80
      when "100000111011" =>  data <= "10100010";  -- 83B = A2
      when "100000111100" =>  data <= "00000000";  -- 83C = 0
      when "100000111101" =>  data <= "11101000";  -- 83D = E8
      when "100000111110" =>  data <= "11101000";  -- 83E = E8
      when "100000111111" =>  data <= "11101000";  -- 83F = E8
      when "100001000000" =>  data <= "11101000";  -- 840 = E8
      when "100001000001" =>  data <= "11101000";  -- 841 = E8
      when "100001000010" =>  data <= "11101000";  -- 842 = E8
      when "100001000011" =>  data <= "11101000";  -- 843 = E8
      when "100001000100" =>  data <= "11101000";  -- 844 = E8
      when "100001000101" =>  data <= "11101000";  -- 845 = E8
      when "100001000110" =>  data <= "11101000";  -- 846 = E8
      when "100001000111" =>  data <= "11101000";  -- 847 = E8
      when "100001001000" =>  data <= "11101000";  -- 848 = E8
      when "100001001001" =>  data <= "11101000";  -- 849 = E8
      when "100001001010" =>  data <= "11101000";  -- 84A = E8
      when "100001001011" =>  data <= "11101000";  -- 84B = E8
      when "100001001100" =>  data <= "11101000";  -- 84C = E8
      when "100001001101" =>  data <= "11100000";  -- 84D = E0
      when "100001001110" =>  data <= "00010000";  -- 84E = 10
      when "100001001111" =>  data <= "11110000";  -- 84F = F0
      when "100001010000" =>  data <= "00000101";  -- 850 = 5
      when "100001010001" =>  data <= "10101001";  -- 851 = A9
      when "100001010010" =>  data <= "01100100";  -- 852 = 64
      when "100001010011" =>  data <= "01001100";  -- 853 = 4C
      when "100001010100" =>  data <= "01000001";  -- 854 = 41
      when "100001010101" =>  data <= "11111001";  -- 855 = F9
      when "100001010110" =>  data <= "10100101";  -- 856 = A5
      when "100001010111" =>  data <= "00000111";  -- 857 = 7
      when "100001011000" =>  data <= "11001001";  -- 858 = C9
      when "100001011001" =>  data <= "00000001";  -- 859 = 1
      when "100001011010" =>  data <= "11110000";  -- 85A = F0
      when "100001011011" =>  data <= "00000101";  -- 85B = 5
      when "100001011100" =>  data <= "10101001";  -- 85C = A9
      when "100001011101" =>  data <= "01100101";  -- 85D = 65
      when "100001011110" =>  data <= "01001100";  -- 85E = 4C
      when "100001011111" =>  data <= "01000001";  -- 85F = 41
      when "100001100000" =>  data <= "11111001";  -- 860 = F9
      when "100001100001" =>  data <= "10101001";  -- 861 = A9
      when "100001100010" =>  data <= "00000000";  -- 862 = 0
      when "100001100011" =>  data <= "10000101";  -- 863 = 85
      when "100001100100" =>  data <= "00000110";  -- 864 = 6
      when "100001100101" =>  data <= "10001101";  -- 865 = 8D
      when "100001100110" =>  data <= "00000111";  -- 866 = 7
      when "100001100111" =>  data <= "10000000";  -- 867 = 80
      when "100001101000" =>  data <= "10101001";  -- 868 = A9
      when "100001101001" =>  data <= "01000100";  -- 869 = 44
      when "100001101010" =>  data <= "10001101";  -- 86A = 8D
      when "100001101011" =>  data <= "00000001";  -- 86B = 1
      when "100001101100" =>  data <= "10000000";  -- 86C = 80
      when "100001101101" =>  data <= "01001100";  -- 86D = 4C
      when "100001101110" =>  data <= "01110011";  -- 86E = 73
      when "100001101111" =>  data <= "11111000";  -- 86F = F8
      when "100001110000" =>  data <= "01001100";  -- 870 = 4C
      when "100001110001" =>  data <= "01111110";  -- 871 = 7E
      when "100001110010" =>  data <= "11111000";  -- 872 = F8
      when "100001110011" =>  data <= "00111000";  -- 873 = 38
      when "100001110100" =>  data <= "10110000";  -- 874 = B0
      when "100001110101" =>  data <= "11111010";  -- 875 = FA
      when "100001110110" =>  data <= "11101010";  -- 876 = EA
      when "100001110111" =>  data <= "11101010";  -- 877 = EA
      when "100001111000" =>  data <= "11101010";  -- 878 = EA
      when "100001111001" =>  data <= "10101001";  -- 879 = A9
      when "100001111010" =>  data <= "01100110";  -- 87A = 66
      when "100001111011" =>  data <= "01001100";  -- 87B = 4C
      when "100001111100" =>  data <= "01000001";  -- 87C = 41
      when "100001111101" =>  data <= "11111001";  -- 87D = F9
      when "100001111110" =>  data <= "10101001";  -- 87E = A9
      when "100001111111" =>  data <= "01000101";  -- 87F = 45
      when "100010000000" =>  data <= "10001101";  -- 880 = 8D
      when "100010000001" =>  data <= "00000001";  -- 881 = 1
      when "100010000010" =>  data <= "10000000";  -- 882 = 80
      when "100010000011" =>  data <= "00111000";  -- 883 = 38
      when "100010000100" =>  data <= "10101001";  -- 884 = A9
      when "100010000101" =>  data <= "00110100";  -- 885 = 34
      when "100010000110" =>  data <= "11101001";  -- 886 = E9
      when "100010000111" =>  data <= "01110101";  -- 887 = 75
      when "100010001000" =>  data <= "10010000";  -- 888 = 90
      when "100010001001" =>  data <= "00000101";  -- 889 = 5
      when "100010001010" =>  data <= "10101001";  -- 88A = A9
      when "100010001011" =>  data <= "01100111";  -- 88B = 67
      when "100010001100" =>  data <= "01001100";  -- 88C = 4C
      when "100010001101" =>  data <= "01000001";  -- 88D = 41
      when "100010001110" =>  data <= "11111001";  -- 88E = F9
      when "100010001111" =>  data <= "10101001";  -- 88F = A9
      when "100010010000" =>  data <= "01000110";  -- 890 = 46
      when "100010010001" =>  data <= "10001101";  -- 891 = 8D
      when "100010010010" =>  data <= "00000001";  -- 892 = 1
      when "100010010011" =>  data <= "10000000";  -- 893 = 80
      when "100010010100" =>  data <= "10111010";  -- 894 = BA
      when "100010010101" =>  data <= "10000110";  -- 895 = 86
      when "100010010110" =>  data <= "00000000";  -- 896 = 0
      when "100010010111" =>  data <= "10101001";  -- 897 = A9
      when "100010011000" =>  data <= "01000010";  -- 898 = 42
      when "100010011001" =>  data <= "01001000";  -- 899 = 48
      when "100010011010" =>  data <= "10101001";  -- 89A = A9
      when "100010011011" =>  data <= "00000000";  -- 89B = 0
      when "100010011100" =>  data <= "10111010";  -- 89C = BA
      when "100010011101" =>  data <= "11101000";  -- 89D = E8
      when "100010011110" =>  data <= "10111101";  -- 89E = BD
      when "100010011111" =>  data <= "00000000";  -- 89F = 0
      when "100010100000" =>  data <= "00000001";  -- 8A0 = 1
      when "100010100001" =>  data <= "11001001";  -- 8A1 = C9
      when "100010100010" =>  data <= "01000010";  -- 8A2 = 42
      when "100010100011" =>  data <= "11110000";  -- 8A3 = F0
      when "100010100100" =>  data <= "00000101";  -- 8A4 = 5
      when "100010100101" =>  data <= "10101001";  -- 8A5 = A9
      when "100010100110" =>  data <= "01101000";  -- 8A6 = 68
      when "100010100111" =>  data <= "01001100";  -- 8A7 = 4C
      when "100010101000" =>  data <= "01000001";  -- 8A8 = 41
      when "100010101001" =>  data <= "11111001";  -- 8A9 = F9
      when "100010101010" =>  data <= "10101001";  -- 8AA = A9
      when "100010101011" =>  data <= "01101001";  -- 8AB = 69
      when "100010101100" =>  data <= "10001101";  -- 8AC = 8D
      when "100010101101" =>  data <= "00010010";  -- 8AD = 12
      when "100010101110" =>  data <= "00000001";  -- 8AE = 1
      when "100010101111" =>  data <= "10101001";  -- 8AF = A9
      when "100010110000" =>  data <= "00000000";  -- 8B0 = 0
      when "100010110001" =>  data <= "10100010";  -- 8B1 = A2
      when "100010110010" =>  data <= "00010001";  -- 8B2 = 11
      when "100010110011" =>  data <= "10011010";  -- 8B3 = 9A
      when "100010110100" =>  data <= "01101000";  -- 8B4 = 68
      when "100010110101" =>  data <= "11001001";  -- 8B5 = C9
      when "100010110110" =>  data <= "01101001";  -- 8B6 = 69
      when "100010110111" =>  data <= "11110000";  -- 8B7 = F0
      when "100010111000" =>  data <= "00000101";  -- 8B8 = 5
      when "100010111001" =>  data <= "10101001";  -- 8B9 = A9
      when "100010111010" =>  data <= "01101001";  -- 8BA = 69
      when "100010111011" =>  data <= "01001100";  -- 8BB = 4C
      when "100010111100" =>  data <= "01000001";  -- 8BC = 41
      when "100010111101" =>  data <= "11111001";  -- 8BD = F9
      when "100010111110" =>  data <= "10100110";  -- 8BE = A6
      when "100010111111" =>  data <= "00000000";  -- 8BF = 0
      when "100011000000" =>  data <= "10011010";  -- 8C0 = 9A
      when "100011000001" =>  data <= "10101001";  -- 8C1 = A9
      when "100011000010" =>  data <= "01000111";  -- 8C2 = 47
      when "100011000011" =>  data <= "10001101";  -- 8C3 = 8D
      when "100011000100" =>  data <= "00000001";  -- 8C4 = 1
      when "100011000101" =>  data <= "10000000";  -- 8C5 = 80
      when "100011000110" =>  data <= "10101001";  -- 8C6 = A9
      when "100011000111" =>  data <= "00000000";  -- 8C7 = 0
      when "100011001000" =>  data <= "01001000";  -- 8C8 = 48
      when "100011001001" =>  data <= "00101000";  -- 8C9 = 28
      when "100011001010" =>  data <= "10000110";  -- 8CA = 86
      when "100011001011" =>  data <= "00001000";  -- 8CB = 8
      when "100011001100" =>  data <= "10101001";  -- 8CC = A9
      when "100011001101" =>  data <= "00000000";  -- 8CD = 0
      when "100011001110" =>  data <= "10000101";  -- 8CE = 85
      when "100011001111" =>  data <= "00000101";  -- 8CF = 5
      when "100011010000" =>  data <= "10101001";  -- 8D0 = A9
      when "100011010001" =>  data <= "00000001";  -- 8D1 = 1
      when "100011010010" =>  data <= "10000101";  -- 8D2 = 85
      when "100011010011" =>  data <= "00000100";  -- 8D3 = 4
      when "100011010100" =>  data <= "10100010";  -- 8D4 = A2
      when "100011010101" =>  data <= "01011001";  -- 8D5 = 59
      when "100011010110" =>  data <= "00000000";  -- 8D6 = 0
      when "100011010111" =>  data <= "11101000";  -- 8D7 = E8
      when "100011011000" =>  data <= "10101001";  -- 8D8 = A9
      when "100011011001" =>  data <= "00000000";  -- 8D9 = 0
      when "100011011010" =>  data <= "10000101";  -- 8DA = 85
      when "100011011011" =>  data <= "00000100";  -- 8DB = 4
      when "100011011100" =>  data <= "10100101";  -- 8DC = A5
      when "100011011101" =>  data <= "00000101";  -- 8DD = 5
      when "100011011110" =>  data <= "11001001";  -- 8DE = C9
      when "100011011111" =>  data <= "00000001";  -- 8DF = 1
      when "100011100000" =>  data <= "11110000";  -- 8E0 = F0
      when "100011100001" =>  data <= "00000101";  -- 8E1 = 5
      when "100011100010" =>  data <= "10101001";  -- 8E2 = A9
      when "100011100011" =>  data <= "01110000";  -- 8E3 = 70
      when "100011100100" =>  data <= "01001100";  -- 8E4 = 4C
      when "100011100101" =>  data <= "01000001";  -- 8E5 = 41
      when "100011100110" =>  data <= "11111001";  -- 8E6 = F9
      when "100011100111" =>  data <= "10100101";  -- 8E7 = A5
      when "100011101000" =>  data <= "00001000";  -- 8E8 = 8
      when "100011101001" =>  data <= "00101001";  -- 8E9 = 29
      when "100011101010" =>  data <= "00010000";  -- 8EA = 10
      when "100011101011" =>  data <= "11010000";  -- 8EB = D0
      when "100011101100" =>  data <= "00000101";  -- 8EC = 5
      when "100011101101" =>  data <= "10101001";  -- 8ED = A9
      when "100011101110" =>  data <= "01110001";  -- 8EE = 71
      when "100011101111" =>  data <= "01001100";  -- 8EF = 4C
      when "100011110000" =>  data <= "01000001";  -- 8F0 = 41
      when "100011110001" =>  data <= "11111001";  -- 8F1 = F9
      when "100011110010" =>  data <= "11100000";  -- 8F2 = E0
      when "100011110011" =>  data <= "01011001";  -- 8F3 = 59
      when "100011110100" =>  data <= "11110000";  -- 8F4 = F0
      when "100011110101" =>  data <= "00000101";  -- 8F5 = 5
      when "100011110110" =>  data <= "10101001";  -- 8F6 = A9
      when "100011110111" =>  data <= "01110010";  -- 8F7 = 72
      when "100011111000" =>  data <= "01001100";  -- 8F8 = 4C
      when "100011111001" =>  data <= "01000001";  -- 8F9 = 41
      when "100011111010" =>  data <= "11111001";  -- 8FA = F9
      when "100011111011" =>  data <= "10101001";  -- 8FB = A9
      when "100011111100" =>  data <= "01001000";  -- 8FC = 48
      when "100011111101" =>  data <= "10001101";  -- 8FD = 8D
      when "100011111110" =>  data <= "00000001";  -- 8FE = 1
      when "100011111111" =>  data <= "10000000";  -- 8FF = 80
      when "100100000000" =>  data <= "10101001";  -- 900 = A9
      when "100100000001" =>  data <= "01010011";  -- 901 = 53
      when "100100000010" =>  data <= "10000101";  -- 902 = 85
      when "100100000011" =>  data <= "00110000";  -- 903 = 30
      when "100100000100" =>  data <= "10101001";  -- 904 = A9
      when "100100000101" =>  data <= "00000000";  -- 905 = 0
      when "100100000110" =>  data <= "10100010";  -- 906 = A2
      when "100100000111" =>  data <= "01000000";  -- 907 = 40
      when "100100001000" =>  data <= "10110101";  -- 908 = B5
      when "100100001001" =>  data <= "11110000";  -- 909 = F0
      when "100100001010" =>  data <= "11001001";  -- 90A = C9
      when "100100001011" =>  data <= "01010011";  -- 90B = 53
      when "100100001100" =>  data <= "11110000";  -- 90C = F0
      when "100100001101" =>  data <= "00000101";  -- 90D = 5
      when "100100001110" =>  data <= "10101001";  -- 90E = A9
      when "100100001111" =>  data <= "01110011";  -- 90F = 73
      when "100100010000" =>  data <= "01001100";  -- 910 = 4C
      when "100100010001" =>  data <= "01000001";  -- 911 = 41
      when "100100010010" =>  data <= "11111001";  -- 912 = F9
      when "100100010011" =>  data <= "10101001";  -- 913 = A9
      when "100100010100" =>  data <= "01001001";  -- 914 = 49
      when "100100010101" =>  data <= "10001101";  -- 915 = 8D
      when "100100010110" =>  data <= "00000001";  -- 916 = 1
      when "100100010111" =>  data <= "10000000";  -- 917 = 80
      when "100100011000" =>  data <= "00011000";  -- 918 = 18
      when "100100011001" =>  data <= "10101001";  -- 919 = A9
      when "100100011010" =>  data <= "11111111";  -- 91A = FF
      when "100100011011" =>  data <= "01101001";  -- 91B = 69
      when "100100011100" =>  data <= "00000001";  -- 91C = 1
      when "100100011101" =>  data <= "10110000";  -- 91D = B0
      when "100100011110" =>  data <= "00000101";  -- 91E = 5
      when "100100011111" =>  data <= "10101001";  -- 91F = A9
      when "100100100000" =>  data <= "01110100";  -- 920 = 74
      when "100100100001" =>  data <= "01001100";  -- 921 = 4C
      when "100100100010" =>  data <= "01000001";  -- 922 = 41
      when "100100100011" =>  data <= "11111001";  -- 923 = F9
      when "100100100100" =>  data <= "10101001";  -- 924 = A9
      when "100100100101" =>  data <= "01001010";  -- 925 = 4A
      when "100100100110" =>  data <= "10001101";  -- 926 = 8D
      when "100100100111" =>  data <= "00000001";  -- 927 = 1
      when "100100101000" =>  data <= "10000000";  -- 928 = 80
      when "100100101001" =>  data <= "00111000";  -- 929 = 38
      when "100100101010" =>  data <= "10101001";  -- 92A = A9
      when "100100101011" =>  data <= "01111111";  -- 92B = 7F
      when "100100101100" =>  data <= "11101001";  -- 92C = E9
      when "100100101101" =>  data <= "01111110";  -- 92D = 7E
      when "100100101110" =>  data <= "01010000";  -- 92E = 50
      when "100100101111" =>  data <= "00000101";  -- 92F = 5
      when "100100110000" =>  data <= "10101001";  -- 930 = A9
      when "100100110001" =>  data <= "01110101";  -- 931 = 75
      when "100100110010" =>  data <= "01001100";  -- 932 = 4C
      when "100100110011" =>  data <= "01000001";  -- 933 = 41
      when "100100110100" =>  data <= "11111001";  -- 934 = F9
      when "100100110101" =>  data <= "01111000";  -- 935 = 78
      when "100100110110" =>  data <= "10101001";  -- 936 = A9
      when "100100110111" =>  data <= "11111111";  -- 937 = FF
      when "100100111000" =>  data <= "10001101";  -- 938 = 8D
      when "100100111001" =>  data <= "00000001";  -- 939 = 1
      when "100100111010" =>  data <= "10000000";  -- 93A = 80
      when "100100111011" =>  data <= "10001101";  -- 93B = 8D
      when "100100111100" =>  data <= "00000000";  -- 93C = 0
      when "100100111101" =>  data <= "10000000";  -- 93D = 80
      when "100100111110" =>  data <= "01001100";  -- 93E = 4C
      when "100100111111" =>  data <= "00110101";  -- 93F = 35
      when "100101000000" =>  data <= "11111001";  -- 940 = F9
      when "100101000001" =>  data <= "01111000";  -- 941 = 78
      when "100101000010" =>  data <= "10001101";  -- 942 = 8D
      when "100101000011" =>  data <= "00000000";  -- 943 = 0
      when "100101000100" =>  data <= "10000000";  -- 944 = 80
      when "100101000101" =>  data <= "01001100";  -- 945 = 4C
      when "100101000110" =>  data <= "01000001";  -- 946 = 41
      when "100101000111" =>  data <= "11111001";  -- 947 = F9
      when "100101001000" =>  data <= "01001000";  -- 948 = 48
      when "100101001001" =>  data <= "10001010";  -- 949 = 8A
      when "100101001010" =>  data <= "01001000";  -- 94A = 48
      when "100101001011" =>  data <= "10011000";  -- 94B = 98
      when "100101001100" =>  data <= "01001000";  -- 94C = 48
      when "100101001101" =>  data <= "10111010";  -- 94D = BA
      when "100101001110" =>  data <= "11101000";  -- 94E = E8
      when "100101001111" =>  data <= "11101000";  -- 94F = E8
      when "100101010000" =>  data <= "11101000";  -- 950 = E8
      when "100101010001" =>  data <= "11101000";  -- 951 = E8
      when "100101010010" =>  data <= "10111101";  -- 952 = BD
      when "100101010011" =>  data <= "00000000";  -- 953 = 0
      when "100101010100" =>  data <= "00000001";  -- 954 = 1
      when "100101010101" =>  data <= "10000101";  -- 955 = 85
      when "100101010110" =>  data <= "00001000";  -- 956 = 8
      when "100101010111" =>  data <= "10100101";  -- 957 = A5
      when "100101011000" =>  data <= "00000100";  -- 958 = 4
      when "100101011001" =>  data <= "11001001";  -- 959 = C9
      when "100101011010" =>  data <= "00000000";  -- 95A = 0
      when "100101011011" =>  data <= "11010000";  -- 95B = D0
      when "100101011100" =>  data <= "00000101";  -- 95C = 5
      when "100101011101" =>  data <= "10101001";  -- 95D = A9
      when "100101011110" =>  data <= "11100000";  -- 95E = E0
      when "100101011111" =>  data <= "01001100";  -- 95F = 4C
      when "100101100000" =>  data <= "01000001";  -- 960 = 41
      when "100101100001" =>  data <= "11111001";  -- 961 = F9
      when "100101100010" =>  data <= "10001101";  -- 962 = 8D
      when "100101100011" =>  data <= "00000101";  -- 963 = 5
      when "100101100100" =>  data <= "10000000";  -- 964 = 80
      when "100101100101" =>  data <= "11100110";  -- 965 = E6
      when "100101100110" =>  data <= "00000101";  -- 966 = 5
      when "100101100111" =>  data <= "01101000";  -- 967 = 68
      when "100101101000" =>  data <= "10101000";  -- 968 = A8
      when "100101101001" =>  data <= "01101000";  -- 969 = 68
      when "100101101010" =>  data <= "10101010";  -- 96A = AA
      when "100101101011" =>  data <= "01101000";  -- 96B = 68
      when "100101101100" =>  data <= "01000000";  -- 96C = 40
      when "100101101101" =>  data <= "01001000";  -- 96D = 48
      when "100101101110" =>  data <= "10001010";  -- 96E = 8A
      when "100101101111" =>  data <= "01001000";  -- 96F = 48
      when "100101110000" =>  data <= "10011000";  -- 970 = 98
      when "100101110001" =>  data <= "01001000";  -- 971 = 48
      when "100101110010" =>  data <= "10100101";  -- 972 = A5
      when "100101110011" =>  data <= "00000110";  -- 973 = 6
      when "100101110100" =>  data <= "11001001";  -- 974 = C9
      when "100101110101" =>  data <= "00000000";  -- 975 = 0
      when "100101110110" =>  data <= "11010000";  -- 976 = D0
      when "100101110111" =>  data <= "00000101";  -- 977 = 5
      when "100101111000" =>  data <= "10101001";  -- 978 = A9
      when "100101111001" =>  data <= "11100000";  -- 979 = E0
      when "100101111010" =>  data <= "01001100";  -- 97A = 4C
      when "100101111011" =>  data <= "01000001";  -- 97B = 41
      when "100101111100" =>  data <= "11111001";  -- 97C = F9
      when "100101111101" =>  data <= "10001101";  -- 97D = 8D
      when "100101111110" =>  data <= "00000111";  -- 97E = 7
      when "100101111111" =>  data <= "10000000";  -- 97F = 80
      when "100110000000" =>  data <= "11100110";  -- 980 = E6
      when "100110000001" =>  data <= "00000111";  -- 981 = 7
      when "100110000010" =>  data <= "01101000";  -- 982 = 68
      when "100110000011" =>  data <= "10101000";  -- 983 = A8
      when "100110000100" =>  data <= "01101000";  -- 984 = 68
      when "100110000101" =>  data <= "10101010";  -- 985 = AA
      when "100110000110" =>  data <= "01101000";  -- 986 = 68
      when "100110000111" =>  data <= "01000000";  -- 987 = 40
      when "100110001000" =>  data <= "01001100";  -- 988 = 4C
      when "100110001001" =>  data <= "01001000";  -- 989 = 48
      when "100110001010" =>  data <= "11111001";  -- 98A = F9
      when "100110001011" =>  data <= "01001100";  -- 98B = 4C
      when "100110001100" =>  data <= "01101101";  -- 98C = 6D
      when "100110001101" =>  data <= "11111001";  -- 98D = F9
      when "100110001110" =>  data <= "11111111";  -- 98E = FF
      when "100110001111" =>  data <= "11111111";  -- 98F = FF
      when "100110010000" =>  data <= "11111111";  -- 990 = FF
      when "100110010001" =>  data <= "11111111";  -- 991 = FF
      when "100110010010" =>  data <= "11111111";  -- 992 = FF
      when "100110010011" =>  data <= "11111111";  -- 993 = FF
      when "100110010100" =>  data <= "11111111";  -- 994 = FF
      when "100110010101" =>  data <= "11111111";  -- 995 = FF
      when "100110010110" =>  data <= "11111111";  -- 996 = FF
      when "100110010111" =>  data <= "11111111";  -- 997 = FF
      when "100110011000" =>  data <= "11111111";  -- 998 = FF
      when "100110011001" =>  data <= "11111111";  -- 999 = FF
      when "100110011010" =>  data <= "11111111";  -- 99A = FF
      when "100110011011" =>  data <= "11111111";  -- 99B = FF
      when "100110011100" =>  data <= "11111111";  -- 99C = FF
      when "100110011101" =>  data <= "11111111";  -- 99D = FF
      when "100110011110" =>  data <= "11111111";  -- 99E = FF
      when "100110011111" =>  data <= "11111111";  -- 99F = FF
      when "100110100000" =>  data <= "11111111";  -- 9A0 = FF
      when "100110100001" =>  data <= "11111111";  -- 9A1 = FF
      when "100110100010" =>  data <= "11111111";  -- 9A2 = FF
      when "100110100011" =>  data <= "11111111";  -- 9A3 = FF
      when "100110100100" =>  data <= "11111111";  -- 9A4 = FF
      when "100110100101" =>  data <= "11111111";  -- 9A5 = FF
      when "100110100110" =>  data <= "11111111";  -- 9A6 = FF
      when "100110100111" =>  data <= "11111111";  -- 9A7 = FF
      when "100110101000" =>  data <= "11111111";  -- 9A8 = FF
      when "100110101001" =>  data <= "11111111";  -- 9A9 = FF
      when "100110101010" =>  data <= "11111111";  -- 9AA = FF
      when "100110101011" =>  data <= "11111111";  -- 9AB = FF
      when "100110101100" =>  data <= "11111111";  -- 9AC = FF
      when "100110101101" =>  data <= "11111111";  -- 9AD = FF
      when "100110101110" =>  data <= "11111111";  -- 9AE = FF
      when "100110101111" =>  data <= "11111111";  -- 9AF = FF
      when "100110110000" =>  data <= "11111111";  -- 9B0 = FF
      when "100110110001" =>  data <= "11111111";  -- 9B1 = FF
      when "100110110010" =>  data <= "11111111";  -- 9B2 = FF
      when "100110110011" =>  data <= "11111111";  -- 9B3 = FF
      when "100110110100" =>  data <= "11111111";  -- 9B4 = FF
      when "100110110101" =>  data <= "11111111";  -- 9B5 = FF
      when "100110110110" =>  data <= "11111111";  -- 9B6 = FF
      when "100110110111" =>  data <= "11111111";  -- 9B7 = FF
      when "100110111000" =>  data <= "11111111";  -- 9B8 = FF
      when "100110111001" =>  data <= "11111111";  -- 9B9 = FF
      when "100110111010" =>  data <= "11111111";  -- 9BA = FF
      when "100110111011" =>  data <= "11111111";  -- 9BB = FF
      when "100110111100" =>  data <= "11111111";  -- 9BC = FF
      when "100110111101" =>  data <= "11111111";  -- 9BD = FF
      when "100110111110" =>  data <= "11111111";  -- 9BE = FF
      when "100110111111" =>  data <= "11111111";  -- 9BF = FF
      when "100111000000" =>  data <= "11111111";  -- 9C0 = FF
      when "100111000001" =>  data <= "11111111";  -- 9C1 = FF
      when "100111000010" =>  data <= "11111111";  -- 9C2 = FF
      when "100111000011" =>  data <= "11111111";  -- 9C3 = FF
      when "100111000100" =>  data <= "11111111";  -- 9C4 = FF
      when "100111000101" =>  data <= "11111111";  -- 9C5 = FF
      when "100111000110" =>  data <= "11111111";  -- 9C6 = FF
      when "100111000111" =>  data <= "11111111";  -- 9C7 = FF
      when "100111001000" =>  data <= "11111111";  -- 9C8 = FF
      when "100111001001" =>  data <= "11111111";  -- 9C9 = FF
      when "100111001010" =>  data <= "11111111";  -- 9CA = FF
      when "100111001011" =>  data <= "11111111";  -- 9CB = FF
      when "100111001100" =>  data <= "11111111";  -- 9CC = FF
      when "100111001101" =>  data <= "11111111";  -- 9CD = FF
      when "100111001110" =>  data <= "11111111";  -- 9CE = FF
      when "100111001111" =>  data <= "11111111";  -- 9CF = FF
      when "100111010000" =>  data <= "11111111";  -- 9D0 = FF
      when "100111010001" =>  data <= "11111111";  -- 9D1 = FF
      when "100111010010" =>  data <= "11111111";  -- 9D2 = FF
      when "100111010011" =>  data <= "11111111";  -- 9D3 = FF
      when "100111010100" =>  data <= "11111111";  -- 9D4 = FF
      when "100111010101" =>  data <= "11111111";  -- 9D5 = FF
      when "100111010110" =>  data <= "11111111";  -- 9D6 = FF
      when "100111010111" =>  data <= "11111111";  -- 9D7 = FF
      when "100111011000" =>  data <= "11111111";  -- 9D8 = FF
      when "100111011001" =>  data <= "11111111";  -- 9D9 = FF
      when "100111011010" =>  data <= "11111111";  -- 9DA = FF
      when "100111011011" =>  data <= "11111111";  -- 9DB = FF
      when "100111011100" =>  data <= "11111111";  -- 9DC = FF
      when "100111011101" =>  data <= "11111111";  -- 9DD = FF
      when "100111011110" =>  data <= "11111111";  -- 9DE = FF
      when "100111011111" =>  data <= "11111111";  -- 9DF = FF
      when "100111100000" =>  data <= "11111111";  -- 9E0 = FF
      when "100111100001" =>  data <= "11111111";  -- 9E1 = FF
      when "100111100010" =>  data <= "11111111";  -- 9E2 = FF
      when "100111100011" =>  data <= "11111111";  -- 9E3 = FF
      when "100111100100" =>  data <= "11111111";  -- 9E4 = FF
      when "100111100101" =>  data <= "11111111";  -- 9E5 = FF
      when "100111100110" =>  data <= "11111111";  -- 9E6 = FF
      when "100111100111" =>  data <= "11111111";  -- 9E7 = FF
      when "100111101000" =>  data <= "11111111";  -- 9E8 = FF
      when "100111101001" =>  data <= "11111111";  -- 9E9 = FF
      when "100111101010" =>  data <= "11111111";  -- 9EA = FF
      when "100111101011" =>  data <= "11111111";  -- 9EB = FF
      when "100111101100" =>  data <= "11111111";  -- 9EC = FF
      when "100111101101" =>  data <= "11111111";  -- 9ED = FF
      when "100111101110" =>  data <= "11111111";  -- 9EE = FF
      when "100111101111" =>  data <= "11111111";  -- 9EF = FF
      when "100111110000" =>  data <= "11111111";  -- 9F0 = FF
      when "100111110001" =>  data <= "11111111";  -- 9F1 = FF
      when "100111110010" =>  data <= "11111111";  -- 9F2 = FF
      when "100111110011" =>  data <= "11111111";  -- 9F3 = FF
      when "100111110100" =>  data <= "11111111";  -- 9F4 = FF
      when "100111110101" =>  data <= "11111111";  -- 9F5 = FF
      when "100111110110" =>  data <= "11111111";  -- 9F6 = FF
      when "100111110111" =>  data <= "11111111";  -- 9F7 = FF
      when "100111111000" =>  data <= "11111111";  -- 9F8 = FF
      when "100111111001" =>  data <= "11111111";  -- 9F9 = FF
      when "100111111010" =>  data <= "11111111";  -- 9FA = FF
      when "100111111011" =>  data <= "11111111";  -- 9FB = FF
      when "100111111100" =>  data <= "11111111";  -- 9FC = FF
      when "100111111101" =>  data <= "11111111";  -- 9FD = FF
      when "100111111110" =>  data <= "11111111";  -- 9FE = FF
      when "100111111111" =>  data <= "11111111";  -- 9FF = FF
      when "101000000000" =>  data <= "11111111";  -- A00 = FF
      when "101000000001" =>  data <= "11111111";  -- A01 = FF
      when "101000000010" =>  data <= "11111111";  -- A02 = FF
      when "101000000011" =>  data <= "11111111";  -- A03 = FF
      when "101000000100" =>  data <= "11111111";  -- A04 = FF
      when "101000000101" =>  data <= "11111111";  -- A05 = FF
      when "101000000110" =>  data <= "11111111";  -- A06 = FF
      when "101000000111" =>  data <= "11111111";  -- A07 = FF
      when "101000001000" =>  data <= "11111111";  -- A08 = FF
      when "101000001001" =>  data <= "11111111";  -- A09 = FF
      when "101000001010" =>  data <= "11111111";  -- A0A = FF
      when "101000001011" =>  data <= "11111111";  -- A0B = FF
      when "101000001100" =>  data <= "11111111";  -- A0C = FF
      when "101000001101" =>  data <= "11111111";  -- A0D = FF
      when "101000001110" =>  data <= "11111111";  -- A0E = FF
      when "101000001111" =>  data <= "11111111";  -- A0F = FF
      when "101000010000" =>  data <= "11111111";  -- A10 = FF
      when "101000010001" =>  data <= "11111111";  -- A11 = FF
      when "101000010010" =>  data <= "11111111";  -- A12 = FF
      when "101000010011" =>  data <= "11111111";  -- A13 = FF
      when "101000010100" =>  data <= "11111111";  -- A14 = FF
      when "101000010101" =>  data <= "11111111";  -- A15 = FF
      when "101000010110" =>  data <= "11111111";  -- A16 = FF
      when "101000010111" =>  data <= "11111111";  -- A17 = FF
      when "101000011000" =>  data <= "11111111";  -- A18 = FF
      when "101000011001" =>  data <= "11111111";  -- A19 = FF
      when "101000011010" =>  data <= "11111111";  -- A1A = FF
      when "101000011011" =>  data <= "11111111";  -- A1B = FF
      when "101000011100" =>  data <= "11111111";  -- A1C = FF
      when "101000011101" =>  data <= "11111111";  -- A1D = FF
      when "101000011110" =>  data <= "11111111";  -- A1E = FF
      when "101000011111" =>  data <= "11111111";  -- A1F = FF
      when "101000100000" =>  data <= "11111111";  -- A20 = FF
      when "101000100001" =>  data <= "11111111";  -- A21 = FF
      when "101000100010" =>  data <= "11111111";  -- A22 = FF
      when "101000100011" =>  data <= "11111111";  -- A23 = FF
      when "101000100100" =>  data <= "11111111";  -- A24 = FF
      when "101000100101" =>  data <= "11111111";  -- A25 = FF
      when "101000100110" =>  data <= "11111111";  -- A26 = FF
      when "101000100111" =>  data <= "11111111";  -- A27 = FF
      when "101000101000" =>  data <= "11111111";  -- A28 = FF
      when "101000101001" =>  data <= "11111111";  -- A29 = FF
      when "101000101010" =>  data <= "11111111";  -- A2A = FF
      when "101000101011" =>  data <= "11111111";  -- A2B = FF
      when "101000101100" =>  data <= "11111111";  -- A2C = FF
      when "101000101101" =>  data <= "11111111";  -- A2D = FF
      when "101000101110" =>  data <= "11111111";  -- A2E = FF
      when "101000101111" =>  data <= "11111111";  -- A2F = FF
      when "101000110000" =>  data <= "11111111";  -- A30 = FF
      when "101000110001" =>  data <= "11111111";  -- A31 = FF
      when "101000110010" =>  data <= "11111111";  -- A32 = FF
      when "101000110011" =>  data <= "11111111";  -- A33 = FF
      when "101000110100" =>  data <= "11111111";  -- A34 = FF
      when "101000110101" =>  data <= "11111111";  -- A35 = FF
      when "101000110110" =>  data <= "11111111";  -- A36 = FF
      when "101000110111" =>  data <= "11111111";  -- A37 = FF
      when "101000111000" =>  data <= "11111111";  -- A38 = FF
      when "101000111001" =>  data <= "11111111";  -- A39 = FF
      when "101000111010" =>  data <= "11111111";  -- A3A = FF
      when "101000111011" =>  data <= "11111111";  -- A3B = FF
      when "101000111100" =>  data <= "11111111";  -- A3C = FF
      when "101000111101" =>  data <= "11111111";  -- A3D = FF
      when "101000111110" =>  data <= "11111111";  -- A3E = FF
      when "101000111111" =>  data <= "11111111";  -- A3F = FF
      when "101001000000" =>  data <= "11111111";  -- A40 = FF
      when "101001000001" =>  data <= "11111111";  -- A41 = FF
      when "101001000010" =>  data <= "11111111";  -- A42 = FF
      when "101001000011" =>  data <= "11111111";  -- A43 = FF
      when "101001000100" =>  data <= "11111111";  -- A44 = FF
      when "101001000101" =>  data <= "11111111";  -- A45 = FF
      when "101001000110" =>  data <= "11111111";  -- A46 = FF
      when "101001000111" =>  data <= "11111111";  -- A47 = FF
      when "101001001000" =>  data <= "11111111";  -- A48 = FF
      when "101001001001" =>  data <= "11111111";  -- A49 = FF
      when "101001001010" =>  data <= "11111111";  -- A4A = FF
      when "101001001011" =>  data <= "11111111";  -- A4B = FF
      when "101001001100" =>  data <= "11111111";  -- A4C = FF
      when "101001001101" =>  data <= "11111111";  -- A4D = FF
      when "101001001110" =>  data <= "11111111";  -- A4E = FF
      when "101001001111" =>  data <= "11111111";  -- A4F = FF
      when "101001010000" =>  data <= "11111111";  -- A50 = FF
      when "101001010001" =>  data <= "11111111";  -- A51 = FF
      when "101001010010" =>  data <= "11111111";  -- A52 = FF
      when "101001010011" =>  data <= "11111111";  -- A53 = FF
      when "101001010100" =>  data <= "11111111";  -- A54 = FF
      when "101001010101" =>  data <= "11111111";  -- A55 = FF
      when "101001010110" =>  data <= "11111111";  -- A56 = FF
      when "101001010111" =>  data <= "11111111";  -- A57 = FF
      when "101001011000" =>  data <= "11111111";  -- A58 = FF
      when "101001011001" =>  data <= "11111111";  -- A59 = FF
      when "101001011010" =>  data <= "11111111";  -- A5A = FF
      when "101001011011" =>  data <= "11111111";  -- A5B = FF
      when "101001011100" =>  data <= "11111111";  -- A5C = FF
      when "101001011101" =>  data <= "11111111";  -- A5D = FF
      when "101001011110" =>  data <= "11111111";  -- A5E = FF
      when "101001011111" =>  data <= "11111111";  -- A5F = FF
      when "101001100000" =>  data <= "11111111";  -- A60 = FF
      when "101001100001" =>  data <= "11111111";  -- A61 = FF
      when "101001100010" =>  data <= "11111111";  -- A62 = FF
      when "101001100011" =>  data <= "11111111";  -- A63 = FF
      when "101001100100" =>  data <= "11111111";  -- A64 = FF
      when "101001100101" =>  data <= "11111111";  -- A65 = FF
      when "101001100110" =>  data <= "11111111";  -- A66 = FF
      when "101001100111" =>  data <= "11111111";  -- A67 = FF
      when "101001101000" =>  data <= "11111111";  -- A68 = FF
      when "101001101001" =>  data <= "11111111";  -- A69 = FF
      when "101001101010" =>  data <= "11111111";  -- A6A = FF
      when "101001101011" =>  data <= "11111111";  -- A6B = FF
      when "101001101100" =>  data <= "11111111";  -- A6C = FF
      when "101001101101" =>  data <= "11111111";  -- A6D = FF
      when "101001101110" =>  data <= "11111111";  -- A6E = FF
      when "101001101111" =>  data <= "11111111";  -- A6F = FF
      when "101001110000" =>  data <= "11111111";  -- A70 = FF
      when "101001110001" =>  data <= "11111111";  -- A71 = FF
      when "101001110010" =>  data <= "11111111";  -- A72 = FF
      when "101001110011" =>  data <= "11111111";  -- A73 = FF
      when "101001110100" =>  data <= "11111111";  -- A74 = FF
      when "101001110101" =>  data <= "11111111";  -- A75 = FF
      when "101001110110" =>  data <= "11111111";  -- A76 = FF
      when "101001110111" =>  data <= "11111111";  -- A77 = FF
      when "101001111000" =>  data <= "11111111";  -- A78 = FF
      when "101001111001" =>  data <= "11111111";  -- A79 = FF
      when "101001111010" =>  data <= "11111111";  -- A7A = FF
      when "101001111011" =>  data <= "11111111";  -- A7B = FF
      when "101001111100" =>  data <= "11111111";  -- A7C = FF
      when "101001111101" =>  data <= "11111111";  -- A7D = FF
      when "101001111110" =>  data <= "11111111";  -- A7E = FF
      when "101001111111" =>  data <= "11111111";  -- A7F = FF
      when "101010000000" =>  data <= "11111111";  -- A80 = FF
      when "101010000001" =>  data <= "11111111";  -- A81 = FF
      when "101010000010" =>  data <= "11111111";  -- A82 = FF
      when "101010000011" =>  data <= "11111111";  -- A83 = FF
      when "101010000100" =>  data <= "11111111";  -- A84 = FF
      when "101010000101" =>  data <= "11111111";  -- A85 = FF
      when "101010000110" =>  data <= "11111111";  -- A86 = FF
      when "101010000111" =>  data <= "11111111";  -- A87 = FF
      when "101010001000" =>  data <= "11111111";  -- A88 = FF
      when "101010001001" =>  data <= "11111111";  -- A89 = FF
      when "101010001010" =>  data <= "11111111";  -- A8A = FF
      when "101010001011" =>  data <= "11111111";  -- A8B = FF
      when "101010001100" =>  data <= "11111111";  -- A8C = FF
      when "101010001101" =>  data <= "11111111";  -- A8D = FF
      when "101010001110" =>  data <= "11111111";  -- A8E = FF
      when "101010001111" =>  data <= "11111111";  -- A8F = FF
      when "101010010000" =>  data <= "11111111";  -- A90 = FF
      when "101010010001" =>  data <= "11111111";  -- A91 = FF
      when "101010010010" =>  data <= "11111111";  -- A92 = FF
      when "101010010011" =>  data <= "11111111";  -- A93 = FF
      when "101010010100" =>  data <= "11111111";  -- A94 = FF
      when "101010010101" =>  data <= "11111111";  -- A95 = FF
      when "101010010110" =>  data <= "11111111";  -- A96 = FF
      when "101010010111" =>  data <= "11111111";  -- A97 = FF
      when "101010011000" =>  data <= "11111111";  -- A98 = FF
      when "101010011001" =>  data <= "11111111";  -- A99 = FF
      when "101010011010" =>  data <= "11111111";  -- A9A = FF
      when "101010011011" =>  data <= "11111111";  -- A9B = FF
      when "101010011100" =>  data <= "11111111";  -- A9C = FF
      when "101010011101" =>  data <= "11111111";  -- A9D = FF
      when "101010011110" =>  data <= "11111111";  -- A9E = FF
      when "101010011111" =>  data <= "11111111";  -- A9F = FF
      when "101010100000" =>  data <= "11111111";  -- AA0 = FF
      when "101010100001" =>  data <= "11111111";  -- AA1 = FF
      when "101010100010" =>  data <= "11111111";  -- AA2 = FF
      when "101010100011" =>  data <= "11111111";  -- AA3 = FF
      when "101010100100" =>  data <= "11111111";  -- AA4 = FF
      when "101010100101" =>  data <= "11111111";  -- AA5 = FF
      when "101010100110" =>  data <= "11111111";  -- AA6 = FF
      when "101010100111" =>  data <= "11111111";  -- AA7 = FF
      when "101010101000" =>  data <= "11111111";  -- AA8 = FF
      when "101010101001" =>  data <= "11111111";  -- AA9 = FF
      when "101010101010" =>  data <= "11111111";  -- AAA = FF
      when "101010101011" =>  data <= "11111111";  -- AAB = FF
      when "101010101100" =>  data <= "11111111";  -- AAC = FF
      when "101010101101" =>  data <= "11111111";  -- AAD = FF
      when "101010101110" =>  data <= "11111111";  -- AAE = FF
      when "101010101111" =>  data <= "11111111";  -- AAF = FF
      when "101010110000" =>  data <= "11111111";  -- AB0 = FF
      when "101010110001" =>  data <= "11111111";  -- AB1 = FF
      when "101010110010" =>  data <= "11111111";  -- AB2 = FF
      when "101010110011" =>  data <= "11111111";  -- AB3 = FF
      when "101010110100" =>  data <= "11111111";  -- AB4 = FF
      when "101010110101" =>  data <= "11111111";  -- AB5 = FF
      when "101010110110" =>  data <= "11111111";  -- AB6 = FF
      when "101010110111" =>  data <= "11111111";  -- AB7 = FF
      when "101010111000" =>  data <= "11111111";  -- AB8 = FF
      when "101010111001" =>  data <= "11111111";  -- AB9 = FF
      when "101010111010" =>  data <= "11111111";  -- ABA = FF
      when "101010111011" =>  data <= "11111111";  -- ABB = FF
      when "101010111100" =>  data <= "11111111";  -- ABC = FF
      when "101010111101" =>  data <= "11111111";  -- ABD = FF
      when "101010111110" =>  data <= "11111111";  -- ABE = FF
      when "101010111111" =>  data <= "11111111";  -- ABF = FF
      when "101011000000" =>  data <= "11111111";  -- AC0 = FF
      when "101011000001" =>  data <= "11111111";  -- AC1 = FF
      when "101011000010" =>  data <= "11111111";  -- AC2 = FF
      when "101011000011" =>  data <= "11111111";  -- AC3 = FF
      when "101011000100" =>  data <= "11111111";  -- AC4 = FF
      when "101011000101" =>  data <= "11111111";  -- AC5 = FF
      when "101011000110" =>  data <= "11111111";  -- AC6 = FF
      when "101011000111" =>  data <= "11111111";  -- AC7 = FF
      when "101011001000" =>  data <= "11111111";  -- AC8 = FF
      when "101011001001" =>  data <= "11111111";  -- AC9 = FF
      when "101011001010" =>  data <= "11111111";  -- ACA = FF
      when "101011001011" =>  data <= "11111111";  -- ACB = FF
      when "101011001100" =>  data <= "11111111";  -- ACC = FF
      when "101011001101" =>  data <= "11111111";  -- ACD = FF
      when "101011001110" =>  data <= "11111111";  -- ACE = FF
      when "101011001111" =>  data <= "11111111";  -- ACF = FF
      when "101011010000" =>  data <= "11111111";  -- AD0 = FF
      when "101011010001" =>  data <= "11111111";  -- AD1 = FF
      when "101011010010" =>  data <= "11111111";  -- AD2 = FF
      when "101011010011" =>  data <= "11111111";  -- AD3 = FF
      when "101011010100" =>  data <= "11111111";  -- AD4 = FF
      when "101011010101" =>  data <= "11111111";  -- AD5 = FF
      when "101011010110" =>  data <= "11111111";  -- AD6 = FF
      when "101011010111" =>  data <= "11111111";  -- AD7 = FF
      when "101011011000" =>  data <= "11111111";  -- AD8 = FF
      when "101011011001" =>  data <= "11111111";  -- AD9 = FF
      when "101011011010" =>  data <= "11111111";  -- ADA = FF
      when "101011011011" =>  data <= "11111111";  -- ADB = FF
      when "101011011100" =>  data <= "11111111";  -- ADC = FF
      when "101011011101" =>  data <= "11111111";  -- ADD = FF
      when "101011011110" =>  data <= "11111111";  -- ADE = FF
      when "101011011111" =>  data <= "11111111";  -- ADF = FF
      when "101011100000" =>  data <= "11111111";  -- AE0 = FF
      when "101011100001" =>  data <= "11111111";  -- AE1 = FF
      when "101011100010" =>  data <= "11111111";  -- AE2 = FF
      when "101011100011" =>  data <= "11111111";  -- AE3 = FF
      when "101011100100" =>  data <= "11111111";  -- AE4 = FF
      when "101011100101" =>  data <= "11111111";  -- AE5 = FF
      when "101011100110" =>  data <= "11111111";  -- AE6 = FF
      when "101011100111" =>  data <= "11111111";  -- AE7 = FF
      when "101011101000" =>  data <= "11111111";  -- AE8 = FF
      when "101011101001" =>  data <= "11111111";  -- AE9 = FF
      when "101011101010" =>  data <= "11111111";  -- AEA = FF
      when "101011101011" =>  data <= "11111111";  -- AEB = FF
      when "101011101100" =>  data <= "11111111";  -- AEC = FF
      when "101011101101" =>  data <= "11111111";  -- AED = FF
      when "101011101110" =>  data <= "11111111";  -- AEE = FF
      when "101011101111" =>  data <= "11111111";  -- AEF = FF
      when "101011110000" =>  data <= "11111111";  -- AF0 = FF
      when "101011110001" =>  data <= "11111111";  -- AF1 = FF
      when "101011110010" =>  data <= "11111111";  -- AF2 = FF
      when "101011110011" =>  data <= "11111111";  -- AF3 = FF
      when "101011110100" =>  data <= "11111111";  -- AF4 = FF
      when "101011110101" =>  data <= "11111111";  -- AF5 = FF
      when "101011110110" =>  data <= "11111111";  -- AF6 = FF
      when "101011110111" =>  data <= "11111111";  -- AF7 = FF
      when "101011111000" =>  data <= "11111111";  -- AF8 = FF
      when "101011111001" =>  data <= "11111111";  -- AF9 = FF
      when "101011111010" =>  data <= "11111111";  -- AFA = FF
      when "101011111011" =>  data <= "11111111";  -- AFB = FF
      when "101011111100" =>  data <= "11111111";  -- AFC = FF
      when "101011111101" =>  data <= "11111111";  -- AFD = FF
      when "101011111110" =>  data <= "11111111";  -- AFE = FF
      when "101011111111" =>  data <= "11111111";  -- AFF = FF
      when "101100000000" =>  data <= "11111111";  -- B00 = FF
      when "101100000001" =>  data <= "11111111";  -- B01 = FF
      when "101100000010" =>  data <= "11111111";  -- B02 = FF
      when "101100000011" =>  data <= "11111111";  -- B03 = FF
      when "101100000100" =>  data <= "11111111";  -- B04 = FF
      when "101100000101" =>  data <= "11111111";  -- B05 = FF
      when "101100000110" =>  data <= "11111111";  -- B06 = FF
      when "101100000111" =>  data <= "11111111";  -- B07 = FF
      when "101100001000" =>  data <= "11111111";  -- B08 = FF
      when "101100001001" =>  data <= "11111111";  -- B09 = FF
      when "101100001010" =>  data <= "11111111";  -- B0A = FF
      when "101100001011" =>  data <= "11111111";  -- B0B = FF
      when "101100001100" =>  data <= "11111111";  -- B0C = FF
      when "101100001101" =>  data <= "11111111";  -- B0D = FF
      when "101100001110" =>  data <= "11111111";  -- B0E = FF
      when "101100001111" =>  data <= "11111111";  -- B0F = FF
      when "101100010000" =>  data <= "11111111";  -- B10 = FF
      when "101100010001" =>  data <= "11111111";  -- B11 = FF
      when "101100010010" =>  data <= "11111111";  -- B12 = FF
      when "101100010011" =>  data <= "11111111";  -- B13 = FF
      when "101100010100" =>  data <= "11111111";  -- B14 = FF
      when "101100010101" =>  data <= "11111111";  -- B15 = FF
      when "101100010110" =>  data <= "11111111";  -- B16 = FF
      when "101100010111" =>  data <= "11111111";  -- B17 = FF
      when "101100011000" =>  data <= "11111111";  -- B18 = FF
      when "101100011001" =>  data <= "11111111";  -- B19 = FF
      when "101100011010" =>  data <= "11111111";  -- B1A = FF
      when "101100011011" =>  data <= "11111111";  -- B1B = FF
      when "101100011100" =>  data <= "11111111";  -- B1C = FF
      when "101100011101" =>  data <= "11111111";  -- B1D = FF
      when "101100011110" =>  data <= "11111111";  -- B1E = FF
      when "101100011111" =>  data <= "11111111";  -- B1F = FF
      when "101100100000" =>  data <= "11111111";  -- B20 = FF
      when "101100100001" =>  data <= "11111111";  -- B21 = FF
      when "101100100010" =>  data <= "11111111";  -- B22 = FF
      when "101100100011" =>  data <= "11111111";  -- B23 = FF
      when "101100100100" =>  data <= "11111111";  -- B24 = FF
      when "101100100101" =>  data <= "11111111";  -- B25 = FF
      when "101100100110" =>  data <= "11111111";  -- B26 = FF
      when "101100100111" =>  data <= "11111111";  -- B27 = FF
      when "101100101000" =>  data <= "11111111";  -- B28 = FF
      when "101100101001" =>  data <= "11111111";  -- B29 = FF
      when "101100101010" =>  data <= "11111111";  -- B2A = FF
      when "101100101011" =>  data <= "11111111";  -- B2B = FF
      when "101100101100" =>  data <= "11111111";  -- B2C = FF
      when "101100101101" =>  data <= "11111111";  -- B2D = FF
      when "101100101110" =>  data <= "11111111";  -- B2E = FF
      when "101100101111" =>  data <= "11111111";  -- B2F = FF
      when "101100110000" =>  data <= "11111111";  -- B30 = FF
      when "101100110001" =>  data <= "11111111";  -- B31 = FF
      when "101100110010" =>  data <= "11111111";  -- B32 = FF
      when "101100110011" =>  data <= "11111111";  -- B33 = FF
      when "101100110100" =>  data <= "11111111";  -- B34 = FF
      when "101100110101" =>  data <= "11111111";  -- B35 = FF
      when "101100110110" =>  data <= "11111111";  -- B36 = FF
      when "101100110111" =>  data <= "11111111";  -- B37 = FF
      when "101100111000" =>  data <= "11111111";  -- B38 = FF
      when "101100111001" =>  data <= "11111111";  -- B39 = FF
      when "101100111010" =>  data <= "11111111";  -- B3A = FF
      when "101100111011" =>  data <= "11111111";  -- B3B = FF
      when "101100111100" =>  data <= "11111111";  -- B3C = FF
      when "101100111101" =>  data <= "11111111";  -- B3D = FF
      when "101100111110" =>  data <= "11111111";  -- B3E = FF
      when "101100111111" =>  data <= "11111111";  -- B3F = FF
      when "101101000000" =>  data <= "11111111";  -- B40 = FF
      when "101101000001" =>  data <= "11111111";  -- B41 = FF
      when "101101000010" =>  data <= "11111111";  -- B42 = FF
      when "101101000011" =>  data <= "11111111";  -- B43 = FF
      when "101101000100" =>  data <= "11111111";  -- B44 = FF
      when "101101000101" =>  data <= "11111111";  -- B45 = FF
      when "101101000110" =>  data <= "11111111";  -- B46 = FF
      when "101101000111" =>  data <= "11111111";  -- B47 = FF
      when "101101001000" =>  data <= "11111111";  -- B48 = FF
      when "101101001001" =>  data <= "11111111";  -- B49 = FF
      when "101101001010" =>  data <= "11111111";  -- B4A = FF
      when "101101001011" =>  data <= "11111111";  -- B4B = FF
      when "101101001100" =>  data <= "11111111";  -- B4C = FF
      when "101101001101" =>  data <= "11111111";  -- B4D = FF
      when "101101001110" =>  data <= "11111111";  -- B4E = FF
      when "101101001111" =>  data <= "11111111";  -- B4F = FF
      when "101101010000" =>  data <= "11111111";  -- B50 = FF
      when "101101010001" =>  data <= "11111111";  -- B51 = FF
      when "101101010010" =>  data <= "11111111";  -- B52 = FF
      when "101101010011" =>  data <= "11111111";  -- B53 = FF
      when "101101010100" =>  data <= "11111111";  -- B54 = FF
      when "101101010101" =>  data <= "11111111";  -- B55 = FF
      when "101101010110" =>  data <= "11111111";  -- B56 = FF
      when "101101010111" =>  data <= "11111111";  -- B57 = FF
      when "101101011000" =>  data <= "11111111";  -- B58 = FF
      when "101101011001" =>  data <= "11111111";  -- B59 = FF
      when "101101011010" =>  data <= "11111111";  -- B5A = FF
      when "101101011011" =>  data <= "11111111";  -- B5B = FF
      when "101101011100" =>  data <= "11111111";  -- B5C = FF
      when "101101011101" =>  data <= "11111111";  -- B5D = FF
      when "101101011110" =>  data <= "11111111";  -- B5E = FF
      when "101101011111" =>  data <= "11111111";  -- B5F = FF
      when "101101100000" =>  data <= "11111111";  -- B60 = FF
      when "101101100001" =>  data <= "11111111";  -- B61 = FF
      when "101101100010" =>  data <= "11111111";  -- B62 = FF
      when "101101100011" =>  data <= "11111111";  -- B63 = FF
      when "101101100100" =>  data <= "11111111";  -- B64 = FF
      when "101101100101" =>  data <= "11111111";  -- B65 = FF
      when "101101100110" =>  data <= "11111111";  -- B66 = FF
      when "101101100111" =>  data <= "11111111";  -- B67 = FF
      when "101101101000" =>  data <= "11111111";  -- B68 = FF
      when "101101101001" =>  data <= "11111111";  -- B69 = FF
      when "101101101010" =>  data <= "11111111";  -- B6A = FF
      when "101101101011" =>  data <= "11111111";  -- B6B = FF
      when "101101101100" =>  data <= "11111111";  -- B6C = FF
      when "101101101101" =>  data <= "11111111";  -- B6D = FF
      when "101101101110" =>  data <= "11111111";  -- B6E = FF
      when "101101101111" =>  data <= "11111111";  -- B6F = FF
      when "101101110000" =>  data <= "11111111";  -- B70 = FF
      when "101101110001" =>  data <= "11111111";  -- B71 = FF
      when "101101110010" =>  data <= "11111111";  -- B72 = FF
      when "101101110011" =>  data <= "11111111";  -- B73 = FF
      when "101101110100" =>  data <= "11111111";  -- B74 = FF
      when "101101110101" =>  data <= "11111111";  -- B75 = FF
      when "101101110110" =>  data <= "11111111";  -- B76 = FF
      when "101101110111" =>  data <= "11111111";  -- B77 = FF
      when "101101111000" =>  data <= "11111111";  -- B78 = FF
      when "101101111001" =>  data <= "11111111";  -- B79 = FF
      when "101101111010" =>  data <= "11111111";  -- B7A = FF
      when "101101111011" =>  data <= "11111111";  -- B7B = FF
      when "101101111100" =>  data <= "11111111";  -- B7C = FF
      when "101101111101" =>  data <= "11111111";  -- B7D = FF
      when "101101111110" =>  data <= "11111111";  -- B7E = FF
      when "101101111111" =>  data <= "11111111";  -- B7F = FF
      when "101110000000" =>  data <= "11111111";  -- B80 = FF
      when "101110000001" =>  data <= "11111111";  -- B81 = FF
      when "101110000010" =>  data <= "11111111";  -- B82 = FF
      when "101110000011" =>  data <= "11111111";  -- B83 = FF
      when "101110000100" =>  data <= "11111111";  -- B84 = FF
      when "101110000101" =>  data <= "11111111";  -- B85 = FF
      when "101110000110" =>  data <= "11111111";  -- B86 = FF
      when "101110000111" =>  data <= "11111111";  -- B87 = FF
      when "101110001000" =>  data <= "11111111";  -- B88 = FF
      when "101110001001" =>  data <= "11111111";  -- B89 = FF
      when "101110001010" =>  data <= "11111111";  -- B8A = FF
      when "101110001011" =>  data <= "11111111";  -- B8B = FF
      when "101110001100" =>  data <= "11111111";  -- B8C = FF
      when "101110001101" =>  data <= "11111111";  -- B8D = FF
      when "101110001110" =>  data <= "11111111";  -- B8E = FF
      when "101110001111" =>  data <= "11111111";  -- B8F = FF
      when "101110010000" =>  data <= "11111111";  -- B90 = FF
      when "101110010001" =>  data <= "11111111";  -- B91 = FF
      when "101110010010" =>  data <= "11111111";  -- B92 = FF
      when "101110010011" =>  data <= "11111111";  -- B93 = FF
      when "101110010100" =>  data <= "11111111";  -- B94 = FF
      when "101110010101" =>  data <= "11111111";  -- B95 = FF
      when "101110010110" =>  data <= "11111111";  -- B96 = FF
      when "101110010111" =>  data <= "11111111";  -- B97 = FF
      when "101110011000" =>  data <= "11111111";  -- B98 = FF
      when "101110011001" =>  data <= "11111111";  -- B99 = FF
      when "101110011010" =>  data <= "11111111";  -- B9A = FF
      when "101110011011" =>  data <= "11111111";  -- B9B = FF
      when "101110011100" =>  data <= "11111111";  -- B9C = FF
      when "101110011101" =>  data <= "11111111";  -- B9D = FF
      when "101110011110" =>  data <= "11111111";  -- B9E = FF
      when "101110011111" =>  data <= "11111111";  -- B9F = FF
      when "101110100000" =>  data <= "11111111";  -- BA0 = FF
      when "101110100001" =>  data <= "11111111";  -- BA1 = FF
      when "101110100010" =>  data <= "11111111";  -- BA2 = FF
      when "101110100011" =>  data <= "11111111";  -- BA3 = FF
      when "101110100100" =>  data <= "11111111";  -- BA4 = FF
      when "101110100101" =>  data <= "11111111";  -- BA5 = FF
      when "101110100110" =>  data <= "11111111";  -- BA6 = FF
      when "101110100111" =>  data <= "11111111";  -- BA7 = FF
      when "101110101000" =>  data <= "11111111";  -- BA8 = FF
      when "101110101001" =>  data <= "11111111";  -- BA9 = FF
      when "101110101010" =>  data <= "11111111";  -- BAA = FF
      when "101110101011" =>  data <= "11111111";  -- BAB = FF
      when "101110101100" =>  data <= "11111111";  -- BAC = FF
      when "101110101101" =>  data <= "11111111";  -- BAD = FF
      when "101110101110" =>  data <= "11111111";  -- BAE = FF
      when "101110101111" =>  data <= "11111111";  -- BAF = FF
      when "101110110000" =>  data <= "11111111";  -- BB0 = FF
      when "101110110001" =>  data <= "11111111";  -- BB1 = FF
      when "101110110010" =>  data <= "11111111";  -- BB2 = FF
      when "101110110011" =>  data <= "11111111";  -- BB3 = FF
      when "101110110100" =>  data <= "11111111";  -- BB4 = FF
      when "101110110101" =>  data <= "11111111";  -- BB5 = FF
      when "101110110110" =>  data <= "11111111";  -- BB6 = FF
      when "101110110111" =>  data <= "11111111";  -- BB7 = FF
      when "101110111000" =>  data <= "11111111";  -- BB8 = FF
      when "101110111001" =>  data <= "11111111";  -- BB9 = FF
      when "101110111010" =>  data <= "11111111";  -- BBA = FF
      when "101110111011" =>  data <= "11111111";  -- BBB = FF
      when "101110111100" =>  data <= "11111111";  -- BBC = FF
      when "101110111101" =>  data <= "11111111";  -- BBD = FF
      when "101110111110" =>  data <= "11111111";  -- BBE = FF
      when "101110111111" =>  data <= "11111111";  -- BBF = FF
      when "101111000000" =>  data <= "11111111";  -- BC0 = FF
      when "101111000001" =>  data <= "11111111";  -- BC1 = FF
      when "101111000010" =>  data <= "11111111";  -- BC2 = FF
      when "101111000011" =>  data <= "11111111";  -- BC3 = FF
      when "101111000100" =>  data <= "11111111";  -- BC4 = FF
      when "101111000101" =>  data <= "11111111";  -- BC5 = FF
      when "101111000110" =>  data <= "11111111";  -- BC6 = FF
      when "101111000111" =>  data <= "11111111";  -- BC7 = FF
      when "101111001000" =>  data <= "11111111";  -- BC8 = FF
      when "101111001001" =>  data <= "11111111";  -- BC9 = FF
      when "101111001010" =>  data <= "11111111";  -- BCA = FF
      when "101111001011" =>  data <= "11111111";  -- BCB = FF
      when "101111001100" =>  data <= "11111111";  -- BCC = FF
      when "101111001101" =>  data <= "11111111";  -- BCD = FF
      when "101111001110" =>  data <= "11111111";  -- BCE = FF
      when "101111001111" =>  data <= "11111111";  -- BCF = FF
      when "101111010000" =>  data <= "11111111";  -- BD0 = FF
      when "101111010001" =>  data <= "11111111";  -- BD1 = FF
      when "101111010010" =>  data <= "11111111";  -- BD2 = FF
      when "101111010011" =>  data <= "11111111";  -- BD3 = FF
      when "101111010100" =>  data <= "11111111";  -- BD4 = FF
      when "101111010101" =>  data <= "11111111";  -- BD5 = FF
      when "101111010110" =>  data <= "11111111";  -- BD6 = FF
      when "101111010111" =>  data <= "11111111";  -- BD7 = FF
      when "101111011000" =>  data <= "11111111";  -- BD8 = FF
      when "101111011001" =>  data <= "11111111";  -- BD9 = FF
      when "101111011010" =>  data <= "11111111";  -- BDA = FF
      when "101111011011" =>  data <= "11111111";  -- BDB = FF
      when "101111011100" =>  data <= "11111111";  -- BDC = FF
      when "101111011101" =>  data <= "11111111";  -- BDD = FF
      when "101111011110" =>  data <= "11111111";  -- BDE = FF
      when "101111011111" =>  data <= "11111111";  -- BDF = FF
      when "101111100000" =>  data <= "11111111";  -- BE0 = FF
      when "101111100001" =>  data <= "11111111";  -- BE1 = FF
      when "101111100010" =>  data <= "11111111";  -- BE2 = FF
      when "101111100011" =>  data <= "11111111";  -- BE3 = FF
      when "101111100100" =>  data <= "11111111";  -- BE4 = FF
      when "101111100101" =>  data <= "11111111";  -- BE5 = FF
      when "101111100110" =>  data <= "11111111";  -- BE6 = FF
      when "101111100111" =>  data <= "11111111";  -- BE7 = FF
      when "101111101000" =>  data <= "11111111";  -- BE8 = FF
      when "101111101001" =>  data <= "11111111";  -- BE9 = FF
      when "101111101010" =>  data <= "11111111";  -- BEA = FF
      when "101111101011" =>  data <= "11111111";  -- BEB = FF
      when "101111101100" =>  data <= "11111111";  -- BEC = FF
      when "101111101101" =>  data <= "11111111";  -- BED = FF
      when "101111101110" =>  data <= "11111111";  -- BEE = FF
      when "101111101111" =>  data <= "11111111";  -- BEF = FF
      when "101111110000" =>  data <= "11111111";  -- BF0 = FF
      when "101111110001" =>  data <= "11111111";  -- BF1 = FF
      when "101111110010" =>  data <= "11111111";  -- BF2 = FF
      when "101111110011" =>  data <= "11111111";  -- BF3 = FF
      when "101111110100" =>  data <= "11111111";  -- BF4 = FF
      when "101111110101" =>  data <= "11111111";  -- BF5 = FF
      when "101111110110" =>  data <= "11111111";  -- BF6 = FF
      when "101111110111" =>  data <= "11111111";  -- BF7 = FF
      when "101111111000" =>  data <= "11111111";  -- BF8 = FF
      when "101111111001" =>  data <= "11111111";  -- BF9 = FF
      when "101111111010" =>  data <= "11111111";  -- BFA = FF
      when "101111111011" =>  data <= "11111111";  -- BFB = FF
      when "101111111100" =>  data <= "11111111";  -- BFC = FF
      when "101111111101" =>  data <= "11111111";  -- BFD = FF
      when "101111111110" =>  data <= "11111111";  -- BFE = FF
      when "101111111111" =>  data <= "11111111";  -- BFF = FF
      when "110000000000" =>  data <= "11111111";  -- C00 = FF
      when "110000000001" =>  data <= "11111111";  -- C01 = FF
      when "110000000010" =>  data <= "11111111";  -- C02 = FF
      when "110000000011" =>  data <= "11111111";  -- C03 = FF
      when "110000000100" =>  data <= "11111111";  -- C04 = FF
      when "110000000101" =>  data <= "11111111";  -- C05 = FF
      when "110000000110" =>  data <= "11111111";  -- C06 = FF
      when "110000000111" =>  data <= "11111111";  -- C07 = FF
      when "110000001000" =>  data <= "11111111";  -- C08 = FF
      when "110000001001" =>  data <= "11111111";  -- C09 = FF
      when "110000001010" =>  data <= "11111111";  -- C0A = FF
      when "110000001011" =>  data <= "11111111";  -- C0B = FF
      when "110000001100" =>  data <= "11111111";  -- C0C = FF
      when "110000001101" =>  data <= "11111111";  -- C0D = FF
      when "110000001110" =>  data <= "11111111";  -- C0E = FF
      when "110000001111" =>  data <= "11111111";  -- C0F = FF
      when "110000010000" =>  data <= "11111111";  -- C10 = FF
      when "110000010001" =>  data <= "11111111";  -- C11 = FF
      when "110000010010" =>  data <= "11111111";  -- C12 = FF
      when "110000010011" =>  data <= "11111111";  -- C13 = FF
      when "110000010100" =>  data <= "11111111";  -- C14 = FF
      when "110000010101" =>  data <= "11111111";  -- C15 = FF
      when "110000010110" =>  data <= "11111111";  -- C16 = FF
      when "110000010111" =>  data <= "11111111";  -- C17 = FF
      when "110000011000" =>  data <= "11111111";  -- C18 = FF
      when "110000011001" =>  data <= "11111111";  -- C19 = FF
      when "110000011010" =>  data <= "11111111";  -- C1A = FF
      when "110000011011" =>  data <= "11111111";  -- C1B = FF
      when "110000011100" =>  data <= "11111111";  -- C1C = FF
      when "110000011101" =>  data <= "11111111";  -- C1D = FF
      when "110000011110" =>  data <= "11111111";  -- C1E = FF
      when "110000011111" =>  data <= "11111111";  -- C1F = FF
      when "110000100000" =>  data <= "11111111";  -- C20 = FF
      when "110000100001" =>  data <= "11111111";  -- C21 = FF
      when "110000100010" =>  data <= "11111111";  -- C22 = FF
      when "110000100011" =>  data <= "11111111";  -- C23 = FF
      when "110000100100" =>  data <= "11111111";  -- C24 = FF
      when "110000100101" =>  data <= "11111111";  -- C25 = FF
      when "110000100110" =>  data <= "11111111";  -- C26 = FF
      when "110000100111" =>  data <= "11111111";  -- C27 = FF
      when "110000101000" =>  data <= "11111111";  -- C28 = FF
      when "110000101001" =>  data <= "11111111";  -- C29 = FF
      when "110000101010" =>  data <= "11111111";  -- C2A = FF
      when "110000101011" =>  data <= "11111111";  -- C2B = FF
      when "110000101100" =>  data <= "11111111";  -- C2C = FF
      when "110000101101" =>  data <= "11111111";  -- C2D = FF
      when "110000101110" =>  data <= "11111111";  -- C2E = FF
      when "110000101111" =>  data <= "11111111";  -- C2F = FF
      when "110000110000" =>  data <= "11111111";  -- C30 = FF
      when "110000110001" =>  data <= "11111111";  -- C31 = FF
      when "110000110010" =>  data <= "11111111";  -- C32 = FF
      when "110000110011" =>  data <= "11111111";  -- C33 = FF
      when "110000110100" =>  data <= "11111111";  -- C34 = FF
      when "110000110101" =>  data <= "11111111";  -- C35 = FF
      when "110000110110" =>  data <= "11111111";  -- C36 = FF
      when "110000110111" =>  data <= "11111111";  -- C37 = FF
      when "110000111000" =>  data <= "11111111";  -- C38 = FF
      when "110000111001" =>  data <= "11111111";  -- C39 = FF
      when "110000111010" =>  data <= "11111111";  -- C3A = FF
      when "110000111011" =>  data <= "11111111";  -- C3B = FF
      when "110000111100" =>  data <= "11111111";  -- C3C = FF
      when "110000111101" =>  data <= "11111111";  -- C3D = FF
      when "110000111110" =>  data <= "11111111";  -- C3E = FF
      when "110000111111" =>  data <= "11111111";  -- C3F = FF
      when "110001000000" =>  data <= "11111111";  -- C40 = FF
      when "110001000001" =>  data <= "11111111";  -- C41 = FF
      when "110001000010" =>  data <= "11111111";  -- C42 = FF
      when "110001000011" =>  data <= "11111111";  -- C43 = FF
      when "110001000100" =>  data <= "11111111";  -- C44 = FF
      when "110001000101" =>  data <= "11111111";  -- C45 = FF
      when "110001000110" =>  data <= "11111111";  -- C46 = FF
      when "110001000111" =>  data <= "11111111";  -- C47 = FF
      when "110001001000" =>  data <= "11111111";  -- C48 = FF
      when "110001001001" =>  data <= "11111111";  -- C49 = FF
      when "110001001010" =>  data <= "11111111";  -- C4A = FF
      when "110001001011" =>  data <= "11111111";  -- C4B = FF
      when "110001001100" =>  data <= "11111111";  -- C4C = FF
      when "110001001101" =>  data <= "11111111";  -- C4D = FF
      when "110001001110" =>  data <= "11111111";  -- C4E = FF
      when "110001001111" =>  data <= "11111111";  -- C4F = FF
      when "110001010000" =>  data <= "11111111";  -- C50 = FF
      when "110001010001" =>  data <= "11111111";  -- C51 = FF
      when "110001010010" =>  data <= "11111111";  -- C52 = FF
      when "110001010011" =>  data <= "11111111";  -- C53 = FF
      when "110001010100" =>  data <= "11111111";  -- C54 = FF
      when "110001010101" =>  data <= "11111111";  -- C55 = FF
      when "110001010110" =>  data <= "11111111";  -- C56 = FF
      when "110001010111" =>  data <= "11111111";  -- C57 = FF
      when "110001011000" =>  data <= "11111111";  -- C58 = FF
      when "110001011001" =>  data <= "11111111";  -- C59 = FF
      when "110001011010" =>  data <= "11111111";  -- C5A = FF
      when "110001011011" =>  data <= "11111111";  -- C5B = FF
      when "110001011100" =>  data <= "11111111";  -- C5C = FF
      when "110001011101" =>  data <= "11111111";  -- C5D = FF
      when "110001011110" =>  data <= "11111111";  -- C5E = FF
      when "110001011111" =>  data <= "11111111";  -- C5F = FF
      when "110001100000" =>  data <= "11111111";  -- C60 = FF
      when "110001100001" =>  data <= "11111111";  -- C61 = FF
      when "110001100010" =>  data <= "11111111";  -- C62 = FF
      when "110001100011" =>  data <= "11111111";  -- C63 = FF
      when "110001100100" =>  data <= "11111111";  -- C64 = FF
      when "110001100101" =>  data <= "11111111";  -- C65 = FF
      when "110001100110" =>  data <= "11111111";  -- C66 = FF
      when "110001100111" =>  data <= "11111111";  -- C67 = FF
      when "110001101000" =>  data <= "11111111";  -- C68 = FF
      when "110001101001" =>  data <= "11111111";  -- C69 = FF
      when "110001101010" =>  data <= "11111111";  -- C6A = FF
      when "110001101011" =>  data <= "11111111";  -- C6B = FF
      when "110001101100" =>  data <= "11111111";  -- C6C = FF
      when "110001101101" =>  data <= "11111111";  -- C6D = FF
      when "110001101110" =>  data <= "11111111";  -- C6E = FF
      when "110001101111" =>  data <= "11111111";  -- C6F = FF
      when "110001110000" =>  data <= "11111111";  -- C70 = FF
      when "110001110001" =>  data <= "11111111";  -- C71 = FF
      when "110001110010" =>  data <= "11111111";  -- C72 = FF
      when "110001110011" =>  data <= "11111111";  -- C73 = FF
      when "110001110100" =>  data <= "11111111";  -- C74 = FF
      when "110001110101" =>  data <= "11111111";  -- C75 = FF
      when "110001110110" =>  data <= "11111111";  -- C76 = FF
      when "110001110111" =>  data <= "11111111";  -- C77 = FF
      when "110001111000" =>  data <= "11111111";  -- C78 = FF
      when "110001111001" =>  data <= "11111111";  -- C79 = FF
      when "110001111010" =>  data <= "11111111";  -- C7A = FF
      when "110001111011" =>  data <= "11111111";  -- C7B = FF
      when "110001111100" =>  data <= "11111111";  -- C7C = FF
      when "110001111101" =>  data <= "11111111";  -- C7D = FF
      when "110001111110" =>  data <= "11111111";  -- C7E = FF
      when "110001111111" =>  data <= "11111111";  -- C7F = FF
      when "110010000000" =>  data <= "11111111";  -- C80 = FF
      when "110010000001" =>  data <= "11111111";  -- C81 = FF
      when "110010000010" =>  data <= "11111111";  -- C82 = FF
      when "110010000011" =>  data <= "11111111";  -- C83 = FF
      when "110010000100" =>  data <= "11111111";  -- C84 = FF
      when "110010000101" =>  data <= "11111111";  -- C85 = FF
      when "110010000110" =>  data <= "11111111";  -- C86 = FF
      when "110010000111" =>  data <= "11111111";  -- C87 = FF
      when "110010001000" =>  data <= "11111111";  -- C88 = FF
      when "110010001001" =>  data <= "11111111";  -- C89 = FF
      when "110010001010" =>  data <= "11111111";  -- C8A = FF
      when "110010001011" =>  data <= "11111111";  -- C8B = FF
      when "110010001100" =>  data <= "11111111";  -- C8C = FF
      when "110010001101" =>  data <= "11111111";  -- C8D = FF
      when "110010001110" =>  data <= "11111111";  -- C8E = FF
      when "110010001111" =>  data <= "11111111";  -- C8F = FF
      when "110010010000" =>  data <= "11111111";  -- C90 = FF
      when "110010010001" =>  data <= "11111111";  -- C91 = FF
      when "110010010010" =>  data <= "11111111";  -- C92 = FF
      when "110010010011" =>  data <= "11111111";  -- C93 = FF
      when "110010010100" =>  data <= "11111111";  -- C94 = FF
      when "110010010101" =>  data <= "11111111";  -- C95 = FF
      when "110010010110" =>  data <= "11111111";  -- C96 = FF
      when "110010010111" =>  data <= "11111111";  -- C97 = FF
      when "110010011000" =>  data <= "11111111";  -- C98 = FF
      when "110010011001" =>  data <= "11111111";  -- C99 = FF
      when "110010011010" =>  data <= "11111111";  -- C9A = FF
      when "110010011011" =>  data <= "11111111";  -- C9B = FF
      when "110010011100" =>  data <= "11111111";  -- C9C = FF
      when "110010011101" =>  data <= "11111111";  -- C9D = FF
      when "110010011110" =>  data <= "11111111";  -- C9E = FF
      when "110010011111" =>  data <= "11111111";  -- C9F = FF
      when "110010100000" =>  data <= "11111111";  -- CA0 = FF
      when "110010100001" =>  data <= "11111111";  -- CA1 = FF
      when "110010100010" =>  data <= "11111111";  -- CA2 = FF
      when "110010100011" =>  data <= "11111111";  -- CA3 = FF
      when "110010100100" =>  data <= "11111111";  -- CA4 = FF
      when "110010100101" =>  data <= "11111111";  -- CA5 = FF
      when "110010100110" =>  data <= "11111111";  -- CA6 = FF
      when "110010100111" =>  data <= "11111111";  -- CA7 = FF
      when "110010101000" =>  data <= "11111111";  -- CA8 = FF
      when "110010101001" =>  data <= "11111111";  -- CA9 = FF
      when "110010101010" =>  data <= "11111111";  -- CAA = FF
      when "110010101011" =>  data <= "11111111";  -- CAB = FF
      when "110010101100" =>  data <= "11111111";  -- CAC = FF
      when "110010101101" =>  data <= "11111111";  -- CAD = FF
      when "110010101110" =>  data <= "11111111";  -- CAE = FF
      when "110010101111" =>  data <= "11111111";  -- CAF = FF
      when "110010110000" =>  data <= "11111111";  -- CB0 = FF
      when "110010110001" =>  data <= "11111111";  -- CB1 = FF
      when "110010110010" =>  data <= "11111111";  -- CB2 = FF
      when "110010110011" =>  data <= "11111111";  -- CB3 = FF
      when "110010110100" =>  data <= "11111111";  -- CB4 = FF
      when "110010110101" =>  data <= "11111111";  -- CB5 = FF
      when "110010110110" =>  data <= "11111111";  -- CB6 = FF
      when "110010110111" =>  data <= "11111111";  -- CB7 = FF
      when "110010111000" =>  data <= "11111111";  -- CB8 = FF
      when "110010111001" =>  data <= "11111111";  -- CB9 = FF
      when "110010111010" =>  data <= "11111111";  -- CBA = FF
      when "110010111011" =>  data <= "11111111";  -- CBB = FF
      when "110010111100" =>  data <= "11111111";  -- CBC = FF
      when "110010111101" =>  data <= "11111111";  -- CBD = FF
      when "110010111110" =>  data <= "11111111";  -- CBE = FF
      when "110010111111" =>  data <= "11111111";  -- CBF = FF
      when "110011000000" =>  data <= "11111111";  -- CC0 = FF
      when "110011000001" =>  data <= "11111111";  -- CC1 = FF
      when "110011000010" =>  data <= "11111111";  -- CC2 = FF
      when "110011000011" =>  data <= "11111111";  -- CC3 = FF
      when "110011000100" =>  data <= "11111111";  -- CC4 = FF
      when "110011000101" =>  data <= "11111111";  -- CC5 = FF
      when "110011000110" =>  data <= "11111111";  -- CC6 = FF
      when "110011000111" =>  data <= "11111111";  -- CC7 = FF
      when "110011001000" =>  data <= "11111111";  -- CC8 = FF
      when "110011001001" =>  data <= "11111111";  -- CC9 = FF
      when "110011001010" =>  data <= "11111111";  -- CCA = FF
      when "110011001011" =>  data <= "11111111";  -- CCB = FF
      when "110011001100" =>  data <= "11111111";  -- CCC = FF
      when "110011001101" =>  data <= "11111111";  -- CCD = FF
      when "110011001110" =>  data <= "11111111";  -- CCE = FF
      when "110011001111" =>  data <= "11111111";  -- CCF = FF
      when "110011010000" =>  data <= "11111111";  -- CD0 = FF
      when "110011010001" =>  data <= "11111111";  -- CD1 = FF
      when "110011010010" =>  data <= "11111111";  -- CD2 = FF
      when "110011010011" =>  data <= "11111111";  -- CD3 = FF
      when "110011010100" =>  data <= "11111111";  -- CD4 = FF
      when "110011010101" =>  data <= "11111111";  -- CD5 = FF
      when "110011010110" =>  data <= "11111111";  -- CD6 = FF
      when "110011010111" =>  data <= "11111111";  -- CD7 = FF
      when "110011011000" =>  data <= "11111111";  -- CD8 = FF
      when "110011011001" =>  data <= "11111111";  -- CD9 = FF
      when "110011011010" =>  data <= "11111111";  -- CDA = FF
      when "110011011011" =>  data <= "11111111";  -- CDB = FF
      when "110011011100" =>  data <= "11111111";  -- CDC = FF
      when "110011011101" =>  data <= "11111111";  -- CDD = FF
      when "110011011110" =>  data <= "11111111";  -- CDE = FF
      when "110011011111" =>  data <= "11111111";  -- CDF = FF
      when "110011100000" =>  data <= "11111111";  -- CE0 = FF
      when "110011100001" =>  data <= "11111111";  -- CE1 = FF
      when "110011100010" =>  data <= "11111111";  -- CE2 = FF
      when "110011100011" =>  data <= "11111111";  -- CE3 = FF
      when "110011100100" =>  data <= "11111111";  -- CE4 = FF
      when "110011100101" =>  data <= "11111111";  -- CE5 = FF
      when "110011100110" =>  data <= "11111111";  -- CE6 = FF
      when "110011100111" =>  data <= "11111111";  -- CE7 = FF
      when "110011101000" =>  data <= "11111111";  -- CE8 = FF
      when "110011101001" =>  data <= "11111111";  -- CE9 = FF
      when "110011101010" =>  data <= "11111111";  -- CEA = FF
      when "110011101011" =>  data <= "11111111";  -- CEB = FF
      when "110011101100" =>  data <= "11111111";  -- CEC = FF
      when "110011101101" =>  data <= "11111111";  -- CED = FF
      when "110011101110" =>  data <= "11111111";  -- CEE = FF
      when "110011101111" =>  data <= "11111111";  -- CEF = FF
      when "110011110000" =>  data <= "11111111";  -- CF0 = FF
      when "110011110001" =>  data <= "11111111";  -- CF1 = FF
      when "110011110010" =>  data <= "11111111";  -- CF2 = FF
      when "110011110011" =>  data <= "11111111";  -- CF3 = FF
      when "110011110100" =>  data <= "11111111";  -- CF4 = FF
      when "110011110101" =>  data <= "11111111";  -- CF5 = FF
      when "110011110110" =>  data <= "11111111";  -- CF6 = FF
      when "110011110111" =>  data <= "11111111";  -- CF7 = FF
      when "110011111000" =>  data <= "11111111";  -- CF8 = FF
      when "110011111001" =>  data <= "11111111";  -- CF9 = FF
      when "110011111010" =>  data <= "11111111";  -- CFA = FF
      when "110011111011" =>  data <= "11111111";  -- CFB = FF
      when "110011111100" =>  data <= "11111111";  -- CFC = FF
      when "110011111101" =>  data <= "11111111";  -- CFD = FF
      when "110011111110" =>  data <= "11111111";  -- CFE = FF
      when "110011111111" =>  data <= "11111111";  -- CFF = FF
      when "110100000000" =>  data <= "11111111";  -- D00 = FF
      when "110100000001" =>  data <= "11111111";  -- D01 = FF
      when "110100000010" =>  data <= "11111111";  -- D02 = FF
      when "110100000011" =>  data <= "11111111";  -- D03 = FF
      when "110100000100" =>  data <= "11111111";  -- D04 = FF
      when "110100000101" =>  data <= "11111111";  -- D05 = FF
      when "110100000110" =>  data <= "11111111";  -- D06 = FF
      when "110100000111" =>  data <= "11111111";  -- D07 = FF
      when "110100001000" =>  data <= "11111111";  -- D08 = FF
      when "110100001001" =>  data <= "11111111";  -- D09 = FF
      when "110100001010" =>  data <= "11111111";  -- D0A = FF
      when "110100001011" =>  data <= "11111111";  -- D0B = FF
      when "110100001100" =>  data <= "11111111";  -- D0C = FF
      when "110100001101" =>  data <= "11111111";  -- D0D = FF
      when "110100001110" =>  data <= "11111111";  -- D0E = FF
      when "110100001111" =>  data <= "11111111";  -- D0F = FF
      when "110100010000" =>  data <= "11111111";  -- D10 = FF
      when "110100010001" =>  data <= "11111111";  -- D11 = FF
      when "110100010010" =>  data <= "11111111";  -- D12 = FF
      when "110100010011" =>  data <= "11111111";  -- D13 = FF
      when "110100010100" =>  data <= "11111111";  -- D14 = FF
      when "110100010101" =>  data <= "11111111";  -- D15 = FF
      when "110100010110" =>  data <= "11111111";  -- D16 = FF
      when "110100010111" =>  data <= "11111111";  -- D17 = FF
      when "110100011000" =>  data <= "11111111";  -- D18 = FF
      when "110100011001" =>  data <= "11111111";  -- D19 = FF
      when "110100011010" =>  data <= "11111111";  -- D1A = FF
      when "110100011011" =>  data <= "11111111";  -- D1B = FF
      when "110100011100" =>  data <= "11111111";  -- D1C = FF
      when "110100011101" =>  data <= "11111111";  -- D1D = FF
      when "110100011110" =>  data <= "11111111";  -- D1E = FF
      when "110100011111" =>  data <= "11111111";  -- D1F = FF
      when "110100100000" =>  data <= "11111111";  -- D20 = FF
      when "110100100001" =>  data <= "11111111";  -- D21 = FF
      when "110100100010" =>  data <= "11111111";  -- D22 = FF
      when "110100100011" =>  data <= "11111111";  -- D23 = FF
      when "110100100100" =>  data <= "11111111";  -- D24 = FF
      when "110100100101" =>  data <= "11111111";  -- D25 = FF
      when "110100100110" =>  data <= "11111111";  -- D26 = FF
      when "110100100111" =>  data <= "11111111";  -- D27 = FF
      when "110100101000" =>  data <= "11111111";  -- D28 = FF
      when "110100101001" =>  data <= "11111111";  -- D29 = FF
      when "110100101010" =>  data <= "11111111";  -- D2A = FF
      when "110100101011" =>  data <= "11111111";  -- D2B = FF
      when "110100101100" =>  data <= "11111111";  -- D2C = FF
      when "110100101101" =>  data <= "11111111";  -- D2D = FF
      when "110100101110" =>  data <= "11111111";  -- D2E = FF
      when "110100101111" =>  data <= "11111111";  -- D2F = FF
      when "110100110000" =>  data <= "11111111";  -- D30 = FF
      when "110100110001" =>  data <= "11111111";  -- D31 = FF
      when "110100110010" =>  data <= "11111111";  -- D32 = FF
      when "110100110011" =>  data <= "11111111";  -- D33 = FF
      when "110100110100" =>  data <= "11111111";  -- D34 = FF
      when "110100110101" =>  data <= "11111111";  -- D35 = FF
      when "110100110110" =>  data <= "11111111";  -- D36 = FF
      when "110100110111" =>  data <= "11111111";  -- D37 = FF
      when "110100111000" =>  data <= "11111111";  -- D38 = FF
      when "110100111001" =>  data <= "11111111";  -- D39 = FF
      when "110100111010" =>  data <= "11111111";  -- D3A = FF
      when "110100111011" =>  data <= "11111111";  -- D3B = FF
      when "110100111100" =>  data <= "11111111";  -- D3C = FF
      when "110100111101" =>  data <= "11111111";  -- D3D = FF
      when "110100111110" =>  data <= "11111111";  -- D3E = FF
      when "110100111111" =>  data <= "11111111";  -- D3F = FF
      when "110101000000" =>  data <= "11111111";  -- D40 = FF
      when "110101000001" =>  data <= "11111111";  -- D41 = FF
      when "110101000010" =>  data <= "11111111";  -- D42 = FF
      when "110101000011" =>  data <= "11111111";  -- D43 = FF
      when "110101000100" =>  data <= "11111111";  -- D44 = FF
      when "110101000101" =>  data <= "11111111";  -- D45 = FF
      when "110101000110" =>  data <= "11111111";  -- D46 = FF
      when "110101000111" =>  data <= "11111111";  -- D47 = FF
      when "110101001000" =>  data <= "11111111";  -- D48 = FF
      when "110101001001" =>  data <= "11111111";  -- D49 = FF
      when "110101001010" =>  data <= "11111111";  -- D4A = FF
      when "110101001011" =>  data <= "11111111";  -- D4B = FF
      when "110101001100" =>  data <= "11111111";  -- D4C = FF
      when "110101001101" =>  data <= "11111111";  -- D4D = FF
      when "110101001110" =>  data <= "11111111";  -- D4E = FF
      when "110101001111" =>  data <= "11111111";  -- D4F = FF
      when "110101010000" =>  data <= "11111111";  -- D50 = FF
      when "110101010001" =>  data <= "11111111";  -- D51 = FF
      when "110101010010" =>  data <= "11111111";  -- D52 = FF
      when "110101010011" =>  data <= "11111111";  -- D53 = FF
      when "110101010100" =>  data <= "11111111";  -- D54 = FF
      when "110101010101" =>  data <= "11111111";  -- D55 = FF
      when "110101010110" =>  data <= "11111111";  -- D56 = FF
      when "110101010111" =>  data <= "11111111";  -- D57 = FF
      when "110101011000" =>  data <= "11111111";  -- D58 = FF
      when "110101011001" =>  data <= "11111111";  -- D59 = FF
      when "110101011010" =>  data <= "11111111";  -- D5A = FF
      when "110101011011" =>  data <= "11111111";  -- D5B = FF
      when "110101011100" =>  data <= "11111111";  -- D5C = FF
      when "110101011101" =>  data <= "11111111";  -- D5D = FF
      when "110101011110" =>  data <= "11111111";  -- D5E = FF
      when "110101011111" =>  data <= "11111111";  -- D5F = FF
      when "110101100000" =>  data <= "11111111";  -- D60 = FF
      when "110101100001" =>  data <= "11111111";  -- D61 = FF
      when "110101100010" =>  data <= "11111111";  -- D62 = FF
      when "110101100011" =>  data <= "11111111";  -- D63 = FF
      when "110101100100" =>  data <= "11111111";  -- D64 = FF
      when "110101100101" =>  data <= "11111111";  -- D65 = FF
      when "110101100110" =>  data <= "11111111";  -- D66 = FF
      when "110101100111" =>  data <= "11111111";  -- D67 = FF
      when "110101101000" =>  data <= "11111111";  -- D68 = FF
      when "110101101001" =>  data <= "11111111";  -- D69 = FF
      when "110101101010" =>  data <= "11111111";  -- D6A = FF
      when "110101101011" =>  data <= "11111111";  -- D6B = FF
      when "110101101100" =>  data <= "11111111";  -- D6C = FF
      when "110101101101" =>  data <= "11111111";  -- D6D = FF
      when "110101101110" =>  data <= "11111111";  -- D6E = FF
      when "110101101111" =>  data <= "11111111";  -- D6F = FF
      when "110101110000" =>  data <= "11111111";  -- D70 = FF
      when "110101110001" =>  data <= "11111111";  -- D71 = FF
      when "110101110010" =>  data <= "11111111";  -- D72 = FF
      when "110101110011" =>  data <= "11111111";  -- D73 = FF
      when "110101110100" =>  data <= "11111111";  -- D74 = FF
      when "110101110101" =>  data <= "11111111";  -- D75 = FF
      when "110101110110" =>  data <= "11111111";  -- D76 = FF
      when "110101110111" =>  data <= "11111111";  -- D77 = FF
      when "110101111000" =>  data <= "11111111";  -- D78 = FF
      when "110101111001" =>  data <= "11111111";  -- D79 = FF
      when "110101111010" =>  data <= "11111111";  -- D7A = FF
      when "110101111011" =>  data <= "11111111";  -- D7B = FF
      when "110101111100" =>  data <= "11111111";  -- D7C = FF
      when "110101111101" =>  data <= "11111111";  -- D7D = FF
      when "110101111110" =>  data <= "11111111";  -- D7E = FF
      when "110101111111" =>  data <= "11111111";  -- D7F = FF
      when "110110000000" =>  data <= "11111111";  -- D80 = FF
      when "110110000001" =>  data <= "11111111";  -- D81 = FF
      when "110110000010" =>  data <= "11111111";  -- D82 = FF
      when "110110000011" =>  data <= "11111111";  -- D83 = FF
      when "110110000100" =>  data <= "11111111";  -- D84 = FF
      when "110110000101" =>  data <= "11111111";  -- D85 = FF
      when "110110000110" =>  data <= "11111111";  -- D86 = FF
      when "110110000111" =>  data <= "11111111";  -- D87 = FF
      when "110110001000" =>  data <= "11111111";  -- D88 = FF
      when "110110001001" =>  data <= "11111111";  -- D89 = FF
      when "110110001010" =>  data <= "11111111";  -- D8A = FF
      when "110110001011" =>  data <= "11111111";  -- D8B = FF
      when "110110001100" =>  data <= "11111111";  -- D8C = FF
      when "110110001101" =>  data <= "11111111";  -- D8D = FF
      when "110110001110" =>  data <= "11111111";  -- D8E = FF
      when "110110001111" =>  data <= "11111111";  -- D8F = FF
      when "110110010000" =>  data <= "11111111";  -- D90 = FF
      when "110110010001" =>  data <= "11111111";  -- D91 = FF
      when "110110010010" =>  data <= "11111111";  -- D92 = FF
      when "110110010011" =>  data <= "11111111";  -- D93 = FF
      when "110110010100" =>  data <= "11111111";  -- D94 = FF
      when "110110010101" =>  data <= "11111111";  -- D95 = FF
      when "110110010110" =>  data <= "11111111";  -- D96 = FF
      when "110110010111" =>  data <= "11111111";  -- D97 = FF
      when "110110011000" =>  data <= "11111111";  -- D98 = FF
      when "110110011001" =>  data <= "11111111";  -- D99 = FF
      when "110110011010" =>  data <= "11111111";  -- D9A = FF
      when "110110011011" =>  data <= "11111111";  -- D9B = FF
      when "110110011100" =>  data <= "11111111";  -- D9C = FF
      when "110110011101" =>  data <= "11111111";  -- D9D = FF
      when "110110011110" =>  data <= "11111111";  -- D9E = FF
      when "110110011111" =>  data <= "11111111";  -- D9F = FF
      when "110110100000" =>  data <= "11111111";  -- DA0 = FF
      when "110110100001" =>  data <= "11111111";  -- DA1 = FF
      when "110110100010" =>  data <= "11111111";  -- DA2 = FF
      when "110110100011" =>  data <= "11111111";  -- DA3 = FF
      when "110110100100" =>  data <= "11111111";  -- DA4 = FF
      when "110110100101" =>  data <= "11111111";  -- DA5 = FF
      when "110110100110" =>  data <= "11111111";  -- DA6 = FF
      when "110110100111" =>  data <= "11111111";  -- DA7 = FF
      when "110110101000" =>  data <= "11111111";  -- DA8 = FF
      when "110110101001" =>  data <= "11111111";  -- DA9 = FF
      when "110110101010" =>  data <= "11111111";  -- DAA = FF
      when "110110101011" =>  data <= "11111111";  -- DAB = FF
      when "110110101100" =>  data <= "11111111";  -- DAC = FF
      when "110110101101" =>  data <= "11111111";  -- DAD = FF
      when "110110101110" =>  data <= "11111111";  -- DAE = FF
      when "110110101111" =>  data <= "11111111";  -- DAF = FF
      when "110110110000" =>  data <= "11111111";  -- DB0 = FF
      when "110110110001" =>  data <= "11111111";  -- DB1 = FF
      when "110110110010" =>  data <= "11111111";  -- DB2 = FF
      when "110110110011" =>  data <= "11111111";  -- DB3 = FF
      when "110110110100" =>  data <= "11111111";  -- DB4 = FF
      when "110110110101" =>  data <= "11111111";  -- DB5 = FF
      when "110110110110" =>  data <= "11111111";  -- DB6 = FF
      when "110110110111" =>  data <= "11111111";  -- DB7 = FF
      when "110110111000" =>  data <= "11111111";  -- DB8 = FF
      when "110110111001" =>  data <= "11111111";  -- DB9 = FF
      when "110110111010" =>  data <= "11111111";  -- DBA = FF
      when "110110111011" =>  data <= "11111111";  -- DBB = FF
      when "110110111100" =>  data <= "11111111";  -- DBC = FF
      when "110110111101" =>  data <= "11111111";  -- DBD = FF
      when "110110111110" =>  data <= "11111111";  -- DBE = FF
      when "110110111111" =>  data <= "11111111";  -- DBF = FF
      when "110111000000" =>  data <= "11111111";  -- DC0 = FF
      when "110111000001" =>  data <= "11111111";  -- DC1 = FF
      when "110111000010" =>  data <= "11111111";  -- DC2 = FF
      when "110111000011" =>  data <= "11111111";  -- DC3 = FF
      when "110111000100" =>  data <= "11111111";  -- DC4 = FF
      when "110111000101" =>  data <= "11111111";  -- DC5 = FF
      when "110111000110" =>  data <= "11111111";  -- DC6 = FF
      when "110111000111" =>  data <= "11111111";  -- DC7 = FF
      when "110111001000" =>  data <= "11111111";  -- DC8 = FF
      when "110111001001" =>  data <= "11111111";  -- DC9 = FF
      when "110111001010" =>  data <= "11111111";  -- DCA = FF
      when "110111001011" =>  data <= "11111111";  -- DCB = FF
      when "110111001100" =>  data <= "11111111";  -- DCC = FF
      when "110111001101" =>  data <= "11111111";  -- DCD = FF
      when "110111001110" =>  data <= "11111111";  -- DCE = FF
      when "110111001111" =>  data <= "11111111";  -- DCF = FF
      when "110111010000" =>  data <= "11111111";  -- DD0 = FF
      when "110111010001" =>  data <= "11111111";  -- DD1 = FF
      when "110111010010" =>  data <= "11111111";  -- DD2 = FF
      when "110111010011" =>  data <= "11111111";  -- DD3 = FF
      when "110111010100" =>  data <= "11111111";  -- DD4 = FF
      when "110111010101" =>  data <= "11111111";  -- DD5 = FF
      when "110111010110" =>  data <= "11111111";  -- DD6 = FF
      when "110111010111" =>  data <= "11111111";  -- DD7 = FF
      when "110111011000" =>  data <= "11111111";  -- DD8 = FF
      when "110111011001" =>  data <= "11111111";  -- DD9 = FF
      when "110111011010" =>  data <= "11111111";  -- DDA = FF
      when "110111011011" =>  data <= "11111111";  -- DDB = FF
      when "110111011100" =>  data <= "11111111";  -- DDC = FF
      when "110111011101" =>  data <= "11111111";  -- DDD = FF
      when "110111011110" =>  data <= "11111111";  -- DDE = FF
      when "110111011111" =>  data <= "11111111";  -- DDF = FF
      when "110111100000" =>  data <= "11111111";  -- DE0 = FF
      when "110111100001" =>  data <= "11111111";  -- DE1 = FF
      when "110111100010" =>  data <= "11111111";  -- DE2 = FF
      when "110111100011" =>  data <= "11111111";  -- DE3 = FF
      when "110111100100" =>  data <= "11111111";  -- DE4 = FF
      when "110111100101" =>  data <= "11111111";  -- DE5 = FF
      when "110111100110" =>  data <= "11111111";  -- DE6 = FF
      when "110111100111" =>  data <= "11111111";  -- DE7 = FF
      when "110111101000" =>  data <= "11111111";  -- DE8 = FF
      when "110111101001" =>  data <= "11111111";  -- DE9 = FF
      when "110111101010" =>  data <= "11111111";  -- DEA = FF
      when "110111101011" =>  data <= "11111111";  -- DEB = FF
      when "110111101100" =>  data <= "11111111";  -- DEC = FF
      when "110111101101" =>  data <= "11111111";  -- DED = FF
      when "110111101110" =>  data <= "11111111";  -- DEE = FF
      when "110111101111" =>  data <= "11111111";  -- DEF = FF
      when "110111110000" =>  data <= "11111111";  -- DF0 = FF
      when "110111110001" =>  data <= "11111111";  -- DF1 = FF
      when "110111110010" =>  data <= "11111111";  -- DF2 = FF
      when "110111110011" =>  data <= "11111111";  -- DF3 = FF
      when "110111110100" =>  data <= "11111111";  -- DF4 = FF
      when "110111110101" =>  data <= "11111111";  -- DF5 = FF
      when "110111110110" =>  data <= "11111111";  -- DF6 = FF
      when "110111110111" =>  data <= "11111111";  -- DF7 = FF
      when "110111111000" =>  data <= "11111111";  -- DF8 = FF
      when "110111111001" =>  data <= "11111111";  -- DF9 = FF
      when "110111111010" =>  data <= "11111111";  -- DFA = FF
      when "110111111011" =>  data <= "11111111";  -- DFB = FF
      when "110111111100" =>  data <= "11111111";  -- DFC = FF
      when "110111111101" =>  data <= "11111111";  -- DFD = FF
      when "110111111110" =>  data <= "11111111";  -- DFE = FF
      when "110111111111" =>  data <= "11111111";  -- DFF = FF
      when "111000000000" =>  data <= "11111111";  -- E00 = FF
      when "111000000001" =>  data <= "11111111";  -- E01 = FF
      when "111000000010" =>  data <= "11111111";  -- E02 = FF
      when "111000000011" =>  data <= "11111111";  -- E03 = FF
      when "111000000100" =>  data <= "11111111";  -- E04 = FF
      when "111000000101" =>  data <= "11111111";  -- E05 = FF
      when "111000000110" =>  data <= "11111111";  -- E06 = FF
      when "111000000111" =>  data <= "11111111";  -- E07 = FF
      when "111000001000" =>  data <= "11111111";  -- E08 = FF
      when "111000001001" =>  data <= "11111111";  -- E09 = FF
      when "111000001010" =>  data <= "11111111";  -- E0A = FF
      when "111000001011" =>  data <= "11111111";  -- E0B = FF
      when "111000001100" =>  data <= "11111111";  -- E0C = FF
      when "111000001101" =>  data <= "11111111";  -- E0D = FF
      when "111000001110" =>  data <= "11111111";  -- E0E = FF
      when "111000001111" =>  data <= "11111111";  -- E0F = FF
      when "111000010000" =>  data <= "11111111";  -- E10 = FF
      when "111000010001" =>  data <= "11111111";  -- E11 = FF
      when "111000010010" =>  data <= "11111111";  -- E12 = FF
      when "111000010011" =>  data <= "11111111";  -- E13 = FF
      when "111000010100" =>  data <= "11111111";  -- E14 = FF
      when "111000010101" =>  data <= "11111111";  -- E15 = FF
      when "111000010110" =>  data <= "11111111";  -- E16 = FF
      when "111000010111" =>  data <= "11111111";  -- E17 = FF
      when "111000011000" =>  data <= "11111111";  -- E18 = FF
      when "111000011001" =>  data <= "11111111";  -- E19 = FF
      when "111000011010" =>  data <= "11111111";  -- E1A = FF
      when "111000011011" =>  data <= "11111111";  -- E1B = FF
      when "111000011100" =>  data <= "11111111";  -- E1C = FF
      when "111000011101" =>  data <= "11111111";  -- E1D = FF
      when "111000011110" =>  data <= "11111111";  -- E1E = FF
      when "111000011111" =>  data <= "11111111";  -- E1F = FF
      when "111000100000" =>  data <= "11111111";  -- E20 = FF
      when "111000100001" =>  data <= "11111111";  -- E21 = FF
      when "111000100010" =>  data <= "11111111";  -- E22 = FF
      when "111000100011" =>  data <= "11111111";  -- E23 = FF
      when "111000100100" =>  data <= "11111111";  -- E24 = FF
      when "111000100101" =>  data <= "11111111";  -- E25 = FF
      when "111000100110" =>  data <= "11111111";  -- E26 = FF
      when "111000100111" =>  data <= "11111111";  -- E27 = FF
      when "111000101000" =>  data <= "11111111";  -- E28 = FF
      when "111000101001" =>  data <= "11111111";  -- E29 = FF
      when "111000101010" =>  data <= "11111111";  -- E2A = FF
      when "111000101011" =>  data <= "11111111";  -- E2B = FF
      when "111000101100" =>  data <= "11111111";  -- E2C = FF
      when "111000101101" =>  data <= "11111111";  -- E2D = FF
      when "111000101110" =>  data <= "11111111";  -- E2E = FF
      when "111000101111" =>  data <= "11111111";  -- E2F = FF
      when "111000110000" =>  data <= "11111111";  -- E30 = FF
      when "111000110001" =>  data <= "11111111";  -- E31 = FF
      when "111000110010" =>  data <= "11111111";  -- E32 = FF
      when "111000110011" =>  data <= "11111111";  -- E33 = FF
      when "111000110100" =>  data <= "11111111";  -- E34 = FF
      when "111000110101" =>  data <= "11111111";  -- E35 = FF
      when "111000110110" =>  data <= "11111111";  -- E36 = FF
      when "111000110111" =>  data <= "11111111";  -- E37 = FF
      when "111000111000" =>  data <= "11111111";  -- E38 = FF
      when "111000111001" =>  data <= "11111111";  -- E39 = FF
      when "111000111010" =>  data <= "11111111";  -- E3A = FF
      when "111000111011" =>  data <= "11111111";  -- E3B = FF
      when "111000111100" =>  data <= "11111111";  -- E3C = FF
      when "111000111101" =>  data <= "11111111";  -- E3D = FF
      when "111000111110" =>  data <= "11111111";  -- E3E = FF
      when "111000111111" =>  data <= "11111111";  -- E3F = FF
      when "111001000000" =>  data <= "11111111";  -- E40 = FF
      when "111001000001" =>  data <= "11111111";  -- E41 = FF
      when "111001000010" =>  data <= "11111111";  -- E42 = FF
      when "111001000011" =>  data <= "11111111";  -- E43 = FF
      when "111001000100" =>  data <= "11111111";  -- E44 = FF
      when "111001000101" =>  data <= "11111111";  -- E45 = FF
      when "111001000110" =>  data <= "11111111";  -- E46 = FF
      when "111001000111" =>  data <= "11111111";  -- E47 = FF
      when "111001001000" =>  data <= "11111111";  -- E48 = FF
      when "111001001001" =>  data <= "11111111";  -- E49 = FF
      when "111001001010" =>  data <= "11111111";  -- E4A = FF
      when "111001001011" =>  data <= "11111111";  -- E4B = FF
      when "111001001100" =>  data <= "11111111";  -- E4C = FF
      when "111001001101" =>  data <= "11111111";  -- E4D = FF
      when "111001001110" =>  data <= "11111111";  -- E4E = FF
      when "111001001111" =>  data <= "11111111";  -- E4F = FF
      when "111001010000" =>  data <= "11111111";  -- E50 = FF
      when "111001010001" =>  data <= "11111111";  -- E51 = FF
      when "111001010010" =>  data <= "11111111";  -- E52 = FF
      when "111001010011" =>  data <= "11111111";  -- E53 = FF
      when "111001010100" =>  data <= "11111111";  -- E54 = FF
      when "111001010101" =>  data <= "11111111";  -- E55 = FF
      when "111001010110" =>  data <= "11111111";  -- E56 = FF
      when "111001010111" =>  data <= "11111111";  -- E57 = FF
      when "111001011000" =>  data <= "11111111";  -- E58 = FF
      when "111001011001" =>  data <= "11111111";  -- E59 = FF
      when "111001011010" =>  data <= "11111111";  -- E5A = FF
      when "111001011011" =>  data <= "11111111";  -- E5B = FF
      when "111001011100" =>  data <= "11111111";  -- E5C = FF
      when "111001011101" =>  data <= "11111111";  -- E5D = FF
      when "111001011110" =>  data <= "11111111";  -- E5E = FF
      when "111001011111" =>  data <= "11111111";  -- E5F = FF
      when "111001100000" =>  data <= "11111111";  -- E60 = FF
      when "111001100001" =>  data <= "11111111";  -- E61 = FF
      when "111001100010" =>  data <= "11111111";  -- E62 = FF
      when "111001100011" =>  data <= "11111111";  -- E63 = FF
      when "111001100100" =>  data <= "11111111";  -- E64 = FF
      when "111001100101" =>  data <= "11111111";  -- E65 = FF
      when "111001100110" =>  data <= "11111111";  -- E66 = FF
      when "111001100111" =>  data <= "11111111";  -- E67 = FF
      when "111001101000" =>  data <= "11111111";  -- E68 = FF
      when "111001101001" =>  data <= "11111111";  -- E69 = FF
      when "111001101010" =>  data <= "11111111";  -- E6A = FF
      when "111001101011" =>  data <= "11111111";  -- E6B = FF
      when "111001101100" =>  data <= "11111111";  -- E6C = FF
      when "111001101101" =>  data <= "11111111";  -- E6D = FF
      when "111001101110" =>  data <= "11111111";  -- E6E = FF
      when "111001101111" =>  data <= "11111111";  -- E6F = FF
      when "111001110000" =>  data <= "11111111";  -- E70 = FF
      when "111001110001" =>  data <= "11111111";  -- E71 = FF
      when "111001110010" =>  data <= "11111111";  -- E72 = FF
      when "111001110011" =>  data <= "11111111";  -- E73 = FF
      when "111001110100" =>  data <= "11111111";  -- E74 = FF
      when "111001110101" =>  data <= "11111111";  -- E75 = FF
      when "111001110110" =>  data <= "11111111";  -- E76 = FF
      when "111001110111" =>  data <= "11111111";  -- E77 = FF
      when "111001111000" =>  data <= "11111111";  -- E78 = FF
      when "111001111001" =>  data <= "11111111";  -- E79 = FF
      when "111001111010" =>  data <= "11111111";  -- E7A = FF
      when "111001111011" =>  data <= "11111111";  -- E7B = FF
      when "111001111100" =>  data <= "11111111";  -- E7C = FF
      when "111001111101" =>  data <= "11111111";  -- E7D = FF
      when "111001111110" =>  data <= "11111111";  -- E7E = FF
      when "111001111111" =>  data <= "11111111";  -- E7F = FF
      when "111010000000" =>  data <= "11111111";  -- E80 = FF
      when "111010000001" =>  data <= "11111111";  -- E81 = FF
      when "111010000010" =>  data <= "11111111";  -- E82 = FF
      when "111010000011" =>  data <= "11111111";  -- E83 = FF
      when "111010000100" =>  data <= "11111111";  -- E84 = FF
      when "111010000101" =>  data <= "11111111";  -- E85 = FF
      when "111010000110" =>  data <= "11111111";  -- E86 = FF
      when "111010000111" =>  data <= "11111111";  -- E87 = FF
      when "111010001000" =>  data <= "11111111";  -- E88 = FF
      when "111010001001" =>  data <= "11111111";  -- E89 = FF
      when "111010001010" =>  data <= "11111111";  -- E8A = FF
      when "111010001011" =>  data <= "11111111";  -- E8B = FF
      when "111010001100" =>  data <= "11111111";  -- E8C = FF
      when "111010001101" =>  data <= "11111111";  -- E8D = FF
      when "111010001110" =>  data <= "11111111";  -- E8E = FF
      when "111010001111" =>  data <= "11111111";  -- E8F = FF
      when "111010010000" =>  data <= "11111111";  -- E90 = FF
      when "111010010001" =>  data <= "11111111";  -- E91 = FF
      when "111010010010" =>  data <= "11111111";  -- E92 = FF
      when "111010010011" =>  data <= "11111111";  -- E93 = FF
      when "111010010100" =>  data <= "11111111";  -- E94 = FF
      when "111010010101" =>  data <= "11111111";  -- E95 = FF
      when "111010010110" =>  data <= "11111111";  -- E96 = FF
      when "111010010111" =>  data <= "11111111";  -- E97 = FF
      when "111010011000" =>  data <= "11111111";  -- E98 = FF
      when "111010011001" =>  data <= "11111111";  -- E99 = FF
      when "111010011010" =>  data <= "11111111";  -- E9A = FF
      when "111010011011" =>  data <= "11111111";  -- E9B = FF
      when "111010011100" =>  data <= "11111111";  -- E9C = FF
      when "111010011101" =>  data <= "11111111";  -- E9D = FF
      when "111010011110" =>  data <= "11111111";  -- E9E = FF
      when "111010011111" =>  data <= "11111111";  -- E9F = FF
      when "111010100000" =>  data <= "11111111";  -- EA0 = FF
      when "111010100001" =>  data <= "11111111";  -- EA1 = FF
      when "111010100010" =>  data <= "11111111";  -- EA2 = FF
      when "111010100011" =>  data <= "11111111";  -- EA3 = FF
      when "111010100100" =>  data <= "11111111";  -- EA4 = FF
      when "111010100101" =>  data <= "11111111";  -- EA5 = FF
      when "111010100110" =>  data <= "11111111";  -- EA6 = FF
      when "111010100111" =>  data <= "11111111";  -- EA7 = FF
      when "111010101000" =>  data <= "11111111";  -- EA8 = FF
      when "111010101001" =>  data <= "11111111";  -- EA9 = FF
      when "111010101010" =>  data <= "11111111";  -- EAA = FF
      when "111010101011" =>  data <= "11111111";  -- EAB = FF
      when "111010101100" =>  data <= "11111111";  -- EAC = FF
      when "111010101101" =>  data <= "11111111";  -- EAD = FF
      when "111010101110" =>  data <= "11111111";  -- EAE = FF
      when "111010101111" =>  data <= "11111111";  -- EAF = FF
      when "111010110000" =>  data <= "11111111";  -- EB0 = FF
      when "111010110001" =>  data <= "11111111";  -- EB1 = FF
      when "111010110010" =>  data <= "11111111";  -- EB2 = FF
      when "111010110011" =>  data <= "11111111";  -- EB3 = FF
      when "111010110100" =>  data <= "11111111";  -- EB4 = FF
      when "111010110101" =>  data <= "11111111";  -- EB5 = FF
      when "111010110110" =>  data <= "11111111";  -- EB6 = FF
      when "111010110111" =>  data <= "11111111";  -- EB7 = FF
      when "111010111000" =>  data <= "11111111";  -- EB8 = FF
      when "111010111001" =>  data <= "11111111";  -- EB9 = FF
      when "111010111010" =>  data <= "11111111";  -- EBA = FF
      when "111010111011" =>  data <= "11111111";  -- EBB = FF
      when "111010111100" =>  data <= "11111111";  -- EBC = FF
      when "111010111101" =>  data <= "11111111";  -- EBD = FF
      when "111010111110" =>  data <= "11111111";  -- EBE = FF
      when "111010111111" =>  data <= "11111111";  -- EBF = FF
      when "111011000000" =>  data <= "11111111";  -- EC0 = FF
      when "111011000001" =>  data <= "11111111";  -- EC1 = FF
      when "111011000010" =>  data <= "11111111";  -- EC2 = FF
      when "111011000011" =>  data <= "11111111";  -- EC3 = FF
      when "111011000100" =>  data <= "11111111";  -- EC4 = FF
      when "111011000101" =>  data <= "11111111";  -- EC5 = FF
      when "111011000110" =>  data <= "11111111";  -- EC6 = FF
      when "111011000111" =>  data <= "11111111";  -- EC7 = FF
      when "111011001000" =>  data <= "11111111";  -- EC8 = FF
      when "111011001001" =>  data <= "11111111";  -- EC9 = FF
      when "111011001010" =>  data <= "11111111";  -- ECA = FF
      when "111011001011" =>  data <= "11111111";  -- ECB = FF
      when "111011001100" =>  data <= "11111111";  -- ECC = FF
      when "111011001101" =>  data <= "11111111";  -- ECD = FF
      when "111011001110" =>  data <= "11111111";  -- ECE = FF
      when "111011001111" =>  data <= "11111111";  -- ECF = FF
      when "111011010000" =>  data <= "11111111";  -- ED0 = FF
      when "111011010001" =>  data <= "11111111";  -- ED1 = FF
      when "111011010010" =>  data <= "11111111";  -- ED2 = FF
      when "111011010011" =>  data <= "11111111";  -- ED3 = FF
      when "111011010100" =>  data <= "11111111";  -- ED4 = FF
      when "111011010101" =>  data <= "11111111";  -- ED5 = FF
      when "111011010110" =>  data <= "11111111";  -- ED6 = FF
      when "111011010111" =>  data <= "11111111";  -- ED7 = FF
      when "111011011000" =>  data <= "11111111";  -- ED8 = FF
      when "111011011001" =>  data <= "11111111";  -- ED9 = FF
      when "111011011010" =>  data <= "11111111";  -- EDA = FF
      when "111011011011" =>  data <= "11111111";  -- EDB = FF
      when "111011011100" =>  data <= "11111111";  -- EDC = FF
      when "111011011101" =>  data <= "11111111";  -- EDD = FF
      when "111011011110" =>  data <= "11111111";  -- EDE = FF
      when "111011011111" =>  data <= "11111111";  -- EDF = FF
      when "111011100000" =>  data <= "11111111";  -- EE0 = FF
      when "111011100001" =>  data <= "11111111";  -- EE1 = FF
      when "111011100010" =>  data <= "11111111";  -- EE2 = FF
      when "111011100011" =>  data <= "11111111";  -- EE3 = FF
      when "111011100100" =>  data <= "11111111";  -- EE4 = FF
      when "111011100101" =>  data <= "11111111";  -- EE5 = FF
      when "111011100110" =>  data <= "11111111";  -- EE6 = FF
      when "111011100111" =>  data <= "11111111";  -- EE7 = FF
      when "111011101000" =>  data <= "11111111";  -- EE8 = FF
      when "111011101001" =>  data <= "11111111";  -- EE9 = FF
      when "111011101010" =>  data <= "11111111";  -- EEA = FF
      when "111011101011" =>  data <= "11111111";  -- EEB = FF
      when "111011101100" =>  data <= "11111111";  -- EEC = FF
      when "111011101101" =>  data <= "11111111";  -- EED = FF
      when "111011101110" =>  data <= "11111111";  -- EEE = FF
      when "111011101111" =>  data <= "11111111";  -- EEF = FF
      when "111011110000" =>  data <= "11111111";  -- EF0 = FF
      when "111011110001" =>  data <= "11111111";  -- EF1 = FF
      when "111011110010" =>  data <= "11111111";  -- EF2 = FF
      when "111011110011" =>  data <= "11111111";  -- EF3 = FF
      when "111011110100" =>  data <= "11111111";  -- EF4 = FF
      when "111011110101" =>  data <= "11111111";  -- EF5 = FF
      when "111011110110" =>  data <= "11111111";  -- EF6 = FF
      when "111011110111" =>  data <= "11111111";  -- EF7 = FF
      when "111011111000" =>  data <= "11111111";  -- EF8 = FF
      when "111011111001" =>  data <= "11111111";  -- EF9 = FF
      when "111011111010" =>  data <= "11111111";  -- EFA = FF
      when "111011111011" =>  data <= "11111111";  -- EFB = FF
      when "111011111100" =>  data <= "11111111";  -- EFC = FF
      when "111011111101" =>  data <= "11111111";  -- EFD = FF
      when "111011111110" =>  data <= "11111111";  -- EFE = FF
      when "111011111111" =>  data <= "11111111";  -- EFF = FF
      when "111100000000" =>  data <= "11111111";  -- F00 = FF
      when "111100000001" =>  data <= "11111111";  -- F01 = FF
      when "111100000010" =>  data <= "11111111";  -- F02 = FF
      when "111100000011" =>  data <= "11111111";  -- F03 = FF
      when "111100000100" =>  data <= "11111111";  -- F04 = FF
      when "111100000101" =>  data <= "11111111";  -- F05 = FF
      when "111100000110" =>  data <= "11111111";  -- F06 = FF
      when "111100000111" =>  data <= "11111111";  -- F07 = FF
      when "111100001000" =>  data <= "11111111";  -- F08 = FF
      when "111100001001" =>  data <= "11111111";  -- F09 = FF
      when "111100001010" =>  data <= "11111111";  -- F0A = FF
      when "111100001011" =>  data <= "11111111";  -- F0B = FF
      when "111100001100" =>  data <= "11111111";  -- F0C = FF
      when "111100001101" =>  data <= "11111111";  -- F0D = FF
      when "111100001110" =>  data <= "11111111";  -- F0E = FF
      when "111100001111" =>  data <= "11111111";  -- F0F = FF
      when "111100010000" =>  data <= "11111111";  -- F10 = FF
      when "111100010001" =>  data <= "11111111";  -- F11 = FF
      when "111100010010" =>  data <= "11111111";  -- F12 = FF
      when "111100010011" =>  data <= "11111111";  -- F13 = FF
      when "111100010100" =>  data <= "11111111";  -- F14 = FF
      when "111100010101" =>  data <= "11111111";  -- F15 = FF
      when "111100010110" =>  data <= "11111111";  -- F16 = FF
      when "111100010111" =>  data <= "11111111";  -- F17 = FF
      when "111100011000" =>  data <= "11111111";  -- F18 = FF
      when "111100011001" =>  data <= "11111111";  -- F19 = FF
      when "111100011010" =>  data <= "11111111";  -- F1A = FF
      when "111100011011" =>  data <= "11111111";  -- F1B = FF
      when "111100011100" =>  data <= "11111111";  -- F1C = FF
      when "111100011101" =>  data <= "11111111";  -- F1D = FF
      when "111100011110" =>  data <= "11111111";  -- F1E = FF
      when "111100011111" =>  data <= "11111111";  -- F1F = FF
      when "111100100000" =>  data <= "11111111";  -- F20 = FF
      when "111100100001" =>  data <= "11111111";  -- F21 = FF
      when "111100100010" =>  data <= "11111111";  -- F22 = FF
      when "111100100011" =>  data <= "11111111";  -- F23 = FF
      when "111100100100" =>  data <= "11111111";  -- F24 = FF
      when "111100100101" =>  data <= "11111111";  -- F25 = FF
      when "111100100110" =>  data <= "11111111";  -- F26 = FF
      when "111100100111" =>  data <= "11111111";  -- F27 = FF
      when "111100101000" =>  data <= "11111111";  -- F28 = FF
      when "111100101001" =>  data <= "11111111";  -- F29 = FF
      when "111100101010" =>  data <= "11111111";  -- F2A = FF
      when "111100101011" =>  data <= "11111111";  -- F2B = FF
      when "111100101100" =>  data <= "11111111";  -- F2C = FF
      when "111100101101" =>  data <= "11111111";  -- F2D = FF
      when "111100101110" =>  data <= "11111111";  -- F2E = FF
      when "111100101111" =>  data <= "11111111";  -- F2F = FF
      when "111100110000" =>  data <= "11111111";  -- F30 = FF
      when "111100110001" =>  data <= "11111111";  -- F31 = FF
      when "111100110010" =>  data <= "11111111";  -- F32 = FF
      when "111100110011" =>  data <= "11111111";  -- F33 = FF
      when "111100110100" =>  data <= "11111111";  -- F34 = FF
      when "111100110101" =>  data <= "11111111";  -- F35 = FF
      when "111100110110" =>  data <= "11111111";  -- F36 = FF
      when "111100110111" =>  data <= "11111111";  -- F37 = FF
      when "111100111000" =>  data <= "11111111";  -- F38 = FF
      when "111100111001" =>  data <= "11111111";  -- F39 = FF
      when "111100111010" =>  data <= "11111111";  -- F3A = FF
      when "111100111011" =>  data <= "11111111";  -- F3B = FF
      when "111100111100" =>  data <= "11111111";  -- F3C = FF
      when "111100111101" =>  data <= "11111111";  -- F3D = FF
      when "111100111110" =>  data <= "11111111";  -- F3E = FF
      when "111100111111" =>  data <= "11111111";  -- F3F = FF
      when "111101000000" =>  data <= "11111111";  -- F40 = FF
      when "111101000001" =>  data <= "11111111";  -- F41 = FF
      when "111101000010" =>  data <= "11111111";  -- F42 = FF
      when "111101000011" =>  data <= "11111111";  -- F43 = FF
      when "111101000100" =>  data <= "11111111";  -- F44 = FF
      when "111101000101" =>  data <= "11111111";  -- F45 = FF
      when "111101000110" =>  data <= "11111111";  -- F46 = FF
      when "111101000111" =>  data <= "11111111";  -- F47 = FF
      when "111101001000" =>  data <= "11111111";  -- F48 = FF
      when "111101001001" =>  data <= "11111111";  -- F49 = FF
      when "111101001010" =>  data <= "11111111";  -- F4A = FF
      when "111101001011" =>  data <= "11111111";  -- F4B = FF
      when "111101001100" =>  data <= "11111111";  -- F4C = FF
      when "111101001101" =>  data <= "11111111";  -- F4D = FF
      when "111101001110" =>  data <= "11111111";  -- F4E = FF
      when "111101001111" =>  data <= "11111111";  -- F4F = FF
      when "111101010000" =>  data <= "11111111";  -- F50 = FF
      when "111101010001" =>  data <= "11111111";  -- F51 = FF
      when "111101010010" =>  data <= "11111111";  -- F52 = FF
      when "111101010011" =>  data <= "11111111";  -- F53 = FF
      when "111101010100" =>  data <= "11111111";  -- F54 = FF
      when "111101010101" =>  data <= "11111111";  -- F55 = FF
      when "111101010110" =>  data <= "11111111";  -- F56 = FF
      when "111101010111" =>  data <= "11111111";  -- F57 = FF
      when "111101011000" =>  data <= "11111111";  -- F58 = FF
      when "111101011001" =>  data <= "11111111";  -- F59 = FF
      when "111101011010" =>  data <= "11111111";  -- F5A = FF
      when "111101011011" =>  data <= "11111111";  -- F5B = FF
      when "111101011100" =>  data <= "11111111";  -- F5C = FF
      when "111101011101" =>  data <= "11111111";  -- F5D = FF
      when "111101011110" =>  data <= "11111111";  -- F5E = FF
      when "111101011111" =>  data <= "11111111";  -- F5F = FF
      when "111101100000" =>  data <= "11111111";  -- F60 = FF
      when "111101100001" =>  data <= "11111111";  -- F61 = FF
      when "111101100010" =>  data <= "11111111";  -- F62 = FF
      when "111101100011" =>  data <= "11111111";  -- F63 = FF
      when "111101100100" =>  data <= "11111111";  -- F64 = FF
      when "111101100101" =>  data <= "11111111";  -- F65 = FF
      when "111101100110" =>  data <= "11111111";  -- F66 = FF
      when "111101100111" =>  data <= "11111111";  -- F67 = FF
      when "111101101000" =>  data <= "11111111";  -- F68 = FF
      when "111101101001" =>  data <= "11111111";  -- F69 = FF
      when "111101101010" =>  data <= "11111111";  -- F6A = FF
      when "111101101011" =>  data <= "11111111";  -- F6B = FF
      when "111101101100" =>  data <= "11111111";  -- F6C = FF
      when "111101101101" =>  data <= "11111111";  -- F6D = FF
      when "111101101110" =>  data <= "11111111";  -- F6E = FF
      when "111101101111" =>  data <= "11111111";  -- F6F = FF
      when "111101110000" =>  data <= "11111111";  -- F70 = FF
      when "111101110001" =>  data <= "11111111";  -- F71 = FF
      when "111101110010" =>  data <= "11111111";  -- F72 = FF
      when "111101110011" =>  data <= "11111111";  -- F73 = FF
      when "111101110100" =>  data <= "11111111";  -- F74 = FF
      when "111101110101" =>  data <= "11111111";  -- F75 = FF
      when "111101110110" =>  data <= "11111111";  -- F76 = FF
      when "111101110111" =>  data <= "11111111";  -- F77 = FF
      when "111101111000" =>  data <= "11111111";  -- F78 = FF
      when "111101111001" =>  data <= "11111111";  -- F79 = FF
      when "111101111010" =>  data <= "11111111";  -- F7A = FF
      when "111101111011" =>  data <= "11111111";  -- F7B = FF
      when "111101111100" =>  data <= "11111111";  -- F7C = FF
      when "111101111101" =>  data <= "11111111";  -- F7D = FF
      when "111101111110" =>  data <= "11111111";  -- F7E = FF
      when "111101111111" =>  data <= "11111111";  -- F7F = FF
      when "111110000000" =>  data <= "11111111";  -- F80 = FF
      when "111110000001" =>  data <= "11111111";  -- F81 = FF
      when "111110000010" =>  data <= "11111111";  -- F82 = FF
      when "111110000011" =>  data <= "11111111";  -- F83 = FF
      when "111110000100" =>  data <= "11111111";  -- F84 = FF
      when "111110000101" =>  data <= "11111111";  -- F85 = FF
      when "111110000110" =>  data <= "11111111";  -- F86 = FF
      when "111110000111" =>  data <= "11111111";  -- F87 = FF
      when "111110001000" =>  data <= "11111111";  -- F88 = FF
      when "111110001001" =>  data <= "11111111";  -- F89 = FF
      when "111110001010" =>  data <= "11111111";  -- F8A = FF
      when "111110001011" =>  data <= "11111111";  -- F8B = FF
      when "111110001100" =>  data <= "11111111";  -- F8C = FF
      when "111110001101" =>  data <= "11111111";  -- F8D = FF
      when "111110001110" =>  data <= "11111111";  -- F8E = FF
      when "111110001111" =>  data <= "11111111";  -- F8F = FF
      when "111110010000" =>  data <= "11111111";  -- F90 = FF
      when "111110010001" =>  data <= "11111111";  -- F91 = FF
      when "111110010010" =>  data <= "11111111";  -- F92 = FF
      when "111110010011" =>  data <= "11111111";  -- F93 = FF
      when "111110010100" =>  data <= "11111111";  -- F94 = FF
      when "111110010101" =>  data <= "11111111";  -- F95 = FF
      when "111110010110" =>  data <= "11111111";  -- F96 = FF
      when "111110010111" =>  data <= "11111111";  -- F97 = FF
      when "111110011000" =>  data <= "11111111";  -- F98 = FF
      when "111110011001" =>  data <= "11111111";  -- F99 = FF
      when "111110011010" =>  data <= "11111111";  -- F9A = FF
      when "111110011011" =>  data <= "11111111";  -- F9B = FF
      when "111110011100" =>  data <= "11111111";  -- F9C = FF
      when "111110011101" =>  data <= "11111111";  -- F9D = FF
      when "111110011110" =>  data <= "11111111";  -- F9E = FF
      when "111110011111" =>  data <= "11111111";  -- F9F = FF
      when "111110100000" =>  data <= "11111111";  -- FA0 = FF
      when "111110100001" =>  data <= "11111111";  -- FA1 = FF
      when "111110100010" =>  data <= "11111111";  -- FA2 = FF
      when "111110100011" =>  data <= "11111111";  -- FA3 = FF
      when "111110100100" =>  data <= "11111111";  -- FA4 = FF
      when "111110100101" =>  data <= "11111111";  -- FA5 = FF
      when "111110100110" =>  data <= "11111111";  -- FA6 = FF
      when "111110100111" =>  data <= "11111111";  -- FA7 = FF
      when "111110101000" =>  data <= "11111111";  -- FA8 = FF
      when "111110101001" =>  data <= "11111111";  -- FA9 = FF
      when "111110101010" =>  data <= "11111111";  -- FAA = FF
      when "111110101011" =>  data <= "11111111";  -- FAB = FF
      when "111110101100" =>  data <= "11111111";  -- FAC = FF
      when "111110101101" =>  data <= "11111111";  -- FAD = FF
      when "111110101110" =>  data <= "11111111";  -- FAE = FF
      when "111110101111" =>  data <= "11111111";  -- FAF = FF
      when "111110110000" =>  data <= "11111111";  -- FB0 = FF
      when "111110110001" =>  data <= "11111111";  -- FB1 = FF
      when "111110110010" =>  data <= "11111111";  -- FB2 = FF
      when "111110110011" =>  data <= "11111111";  -- FB3 = FF
      when "111110110100" =>  data <= "11111111";  -- FB4 = FF
      when "111110110101" =>  data <= "11111111";  -- FB5 = FF
      when "111110110110" =>  data <= "11111111";  -- FB6 = FF
      when "111110110111" =>  data <= "11111111";  -- FB7 = FF
      when "111110111000" =>  data <= "11111111";  -- FB8 = FF
      when "111110111001" =>  data <= "11111111";  -- FB9 = FF
      when "111110111010" =>  data <= "11111111";  -- FBA = FF
      when "111110111011" =>  data <= "11111111";  -- FBB = FF
      when "111110111100" =>  data <= "11111111";  -- FBC = FF
      when "111110111101" =>  data <= "11111111";  -- FBD = FF
      when "111110111110" =>  data <= "11111111";  -- FBE = FF
      when "111110111111" =>  data <= "11111111";  -- FBF = FF
      when "111111000000" =>  data <= "11111111";  -- FC0 = FF
      when "111111000001" =>  data <= "11111111";  -- FC1 = FF
      when "111111000010" =>  data <= "11111111";  -- FC2 = FF
      when "111111000011" =>  data <= "11111111";  -- FC3 = FF
      when "111111000100" =>  data <= "11111111";  -- FC4 = FF
      when "111111000101" =>  data <= "11111111";  -- FC5 = FF
      when "111111000110" =>  data <= "11111111";  -- FC6 = FF
      when "111111000111" =>  data <= "11111111";  -- FC7 = FF
      when "111111001000" =>  data <= "11111111";  -- FC8 = FF
      when "111111001001" =>  data <= "11111111";  -- FC9 = FF
      when "111111001010" =>  data <= "11111111";  -- FCA = FF
      when "111111001011" =>  data <= "11111111";  -- FCB = FF
      when "111111001100" =>  data <= "11111111";  -- FCC = FF
      when "111111001101" =>  data <= "11111111";  -- FCD = FF
      when "111111001110" =>  data <= "11111111";  -- FCE = FF
      when "111111001111" =>  data <= "11111111";  -- FCF = FF
      when "111111010000" =>  data <= "11111111";  -- FD0 = FF
      when "111111010001" =>  data <= "11111111";  -- FD1 = FF
      when "111111010010" =>  data <= "11111111";  -- FD2 = FF
      when "111111010011" =>  data <= "11111111";  -- FD3 = FF
      when "111111010100" =>  data <= "11111111";  -- FD4 = FF
      when "111111010101" =>  data <= "11111111";  -- FD5 = FF
      when "111111010110" =>  data <= "11111111";  -- FD6 = FF
      when "111111010111" =>  data <= "11111111";  -- FD7 = FF
      when "111111011000" =>  data <= "11111111";  -- FD8 = FF
      when "111111011001" =>  data <= "11111111";  -- FD9 = FF
      when "111111011010" =>  data <= "11111111";  -- FDA = FF
      when "111111011011" =>  data <= "11111111";  -- FDB = FF
      when "111111011100" =>  data <= "11111111";  -- FDC = FF
      when "111111011101" =>  data <= "11111111";  -- FDD = FF
      when "111111011110" =>  data <= "11111111";  -- FDE = FF
      when "111111011111" =>  data <= "11111111";  -- FDF = FF
      when "111111100000" =>  data <= "11111111";  -- FE0 = FF
      when "111111100001" =>  data <= "11111111";  -- FE1 = FF
      when "111111100010" =>  data <= "11111111";  -- FE2 = FF
      when "111111100011" =>  data <= "11111111";  -- FE3 = FF
      when "111111100100" =>  data <= "11111111";  -- FE4 = FF
      when "111111100101" =>  data <= "11111111";  -- FE5 = FF
      when "111111100110" =>  data <= "11111111";  -- FE6 = FF
      when "111111100111" =>  data <= "11111111";  -- FE7 = FF
      when "111111101000" =>  data <= "11111111";  -- FE8 = FF
      when "111111101001" =>  data <= "11111111";  -- FE9 = FF
      when "111111101010" =>  data <= "11111111";  -- FEA = FF
      when "111111101011" =>  data <= "11111111";  -- FEB = FF
      when "111111101100" =>  data <= "11111111";  -- FEC = FF
      when "111111101101" =>  data <= "11111111";  -- FED = FF
      when "111111101110" =>  data <= "11111111";  -- FEE = FF
      when "111111101111" =>  data <= "11111111";  -- FEF = FF
      when "111111110000" =>  data <= "11111111";  -- FF0 = FF
      when "111111110001" =>  data <= "11111111";  -- FF1 = FF
      when "111111110010" =>  data <= "11111111";  -- FF2 = FF
      when "111111110011" =>  data <= "11111111";  -- FF3 = FF
      when "111111110100" =>  data <= "11111111";  -- FF4 = FF
      when "111111110101" =>  data <= "11111111";  -- FF5 = FF
      when "111111110110" =>  data <= "11111111";  -- FF6 = FF
      when "111111110111" =>  data <= "11111111";  -- FF7 = FF
      when "111111111000" =>  data <= "11111111";  -- FF8 = FF
      when "111111111001" =>  data <= "11111111";  -- FF9 = FF
      when "111111111010" =>  data <= "10001011";  -- FFA = 8B
      when "111111111011" =>  data <= "11111001";  -- FFB = F9
      when "111111111100" =>  data <= "00000000";  -- FFC = 0
      when "111111111101" =>  data <= "11110000";  -- FFD = F0
      when "111111111110" =>  data <= "10001000";  -- FFE = 88
      when "111111111111" =>  data <= "11111001";  -- FFF = F9
      --end_of_rom
      when others =>  data <= "00000000";
    end case;
  end process;

end arch_test_rom;

------------------------------------------------------------------------------
------------------------------------------------------------------------------

