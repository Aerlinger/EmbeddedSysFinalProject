library ieee;
use ieee.std_l:
