library IEEE;
use IEEE.std_logic_1164.all;

package constants is

	constant Flag_C 	: integer := 0;
	constant Flag_Z 	: integer := 1;
	constant Flag_I 	: integer := 2;
	constant Flag_D 	: integer := 3;
	constant Flag_B 	: integer := 4;
	constant Flag_1 	: integer := 5;
	constant Flag_V 	: integer := 6;
	constant Flag_N 	: integer := 7;

end package;