library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package roms is

	type rom16 	is array (0 to 15) of std_logic_vector(7 downto 0);
	type rom32 	is array (0 to 31) of std_logic_vector(7 downto 0);
	type rom48 	is array (0 to 47) of std_logic_vector(7 downto 0);
	type rom64 	is array (0 to 63) of std_logic_vector(7 downto 0);
	type rom128 is array (0 to 127) of std_logic_vector(7 downto 0);
	type rom256 is array (0 to 255) of std_logic_vector(7 downto 0);
	type rom512 	is array (0 to 15) of std_logic_vector(7 downto 0);
	type rom1024 	is array (0 to 15) of std_logic_vector(7 downto 0);
	
	constant LD_TEST : rom256 :=
	(
		-- the 6 lines below are for the LDA, LDX and LDY opcodes in all the different address modes.
		x"A9", x"11", x"a2", x"22", x"a0", x"33", x"a5", x"20", x"b5", x"20", x"ad", x"21", x"00", x"bd", x"21", x"00",
		x"B9", x"21", x"00", x"a1", x"22", x"b1", x"22", x"ff", x"ff", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"ab", x"33", x"22", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"42", x"43", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"54", x"55", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"66", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --7
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --8
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --9
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --10
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --11
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --12
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --13
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --14
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00" --15
	);
	
	constant INC_DEC_TEST : rom32 := 
	(
		x"EE", x"20", x"00", x"AD", x"20", x"00", x"EE", x"20", x"00", x"AD", x"20", x"00", x"EE", x"20", x"00", x"AD", 
		x"20", x"00", x"CE", x"20", x"00", x"AD", x"20", x"00", x"CE", x"20", x"00", x"AD", x"20", x"00", x"ff", x"ff"
	);
		
	constant CMP_TEST : rom32 := 
	(
		x"EE", x"20", x"00", x"AD", x"20", x"00", x"EE", x"20", x"00", x"AD", x"20", x"00", x"EE", x"20", x"00", x"AD", 
		x"20", x"00", x"CE", x"20", x"00", x"AD", x"20", x"00", x"CE", x"20", x"00", x"AD", x"20", x"00", x"ff", x"ff"
	);
	
	constant JMP_TEST : rom16 := 
	(
		x"ee", x"10", x"00", x"ad", x"10", x"00", x"4c", x"00", x"00", x"ff", x"ff", x"00", x"00", x"00", x"00", x"00"
	);
	
	
	constant BOUNCING_BALL : rom256 :=
	(
		x"A2", x"00", 
		x"A0", x"00", 
		x"A9", x"A0", x"8D", x"70", x"00", 
		x"A9", x"D6", 
		x"8D", x"71", x"00", --Init1/2 (24, x18)
		--		
		x"A9", x"01", x"8D", x"72", x"00", x"A9", x"01", x"8D", x"73", x"00", --Init2/2 (24, x18)
		x"AD", x"72", x"00", x"C9", x"01", x"F0", x"0B", x"D0", x"11", --B1: 0018 (9) --B3 and B4
		x"AD", x"73", x"00", x"C9", x"01", x"F0", x"11", x"D0", x"17", --B2: 0021 (9) --B5 and B6
		x"E8", x"EC", x"70", x"00", 		  x"F0", x"18", x"D0", x"39", --B3: 002A (8) --B7 and B12
		x"CA", x"E0", x"00",               x"F0", x"19", x"D0", x"32", --B4: 0032 (7) --B8 and B120
		x"C8", x"CC", x"71", x"00",        x"F0", x"19", x"D0", x"23", --B5: 0039 (8) --B9 and B11
		x"88", x"C0", x"00",               x"F0", x"1A", x"D0", x"20", --B6: 0041 (7) --B10 and B110
		x"A9", x"00", x"8D", x"72", x"00", x"4C", x"21", x"00", --B7: 0048 (8) --J2
		x"A9", x"01", x"8D", x"72", x"00", x"4C", x"21", x"00", --B8: 0050 (8) --J2
		x"A9", x"00", x"8D", x"73", x"00", x"4C", x"18", x"00", --B9: 0058 (8) --J1
		x"A9", x"01", x"8D", x"73", x"00", x"4C", x"18", x"00", --B10: 0060 (8) --J1
		x"4C", x"18", x"00", --B11: 0068 (3) --J1
		x"4C", x"21", x"00", --B12: 006B (3) --J2
		
		x"ff", x"ff", --6
		
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --7
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --8
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --9
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --10
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --11
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --12
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --13
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", --14
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00" --15
	);
	
end;