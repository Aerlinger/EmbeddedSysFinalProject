------------------------------------------------------------------
---
---  c6502.vhd
---  when         who              what
---  dec12 2003    created         huyvo@comcast.net
---
---
------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity c6502 is

Port (
	clock: in std_logic;
	reset : in std_logic;
	data: inout std_logic_vector(7 downto 0);
	wr:  out std_logic;
	rd: out std_logic;
	ce1: out std_logic;
	
	address: out std_logic_vector(15 downto 0);

-- debug
	--c: out std_logic_vector(3 downto 0)
	peep: out std_logic_vector(7 downto 0)

    );
end c6502;

architecture c6502_architecture of c6502 is


	component IBUFG
		port (
			I : in STD_LOGIC; 
			O : out std_logic
		);
	end component;
 
	------------------------------------------------------------------------
	-- Signal Declarations
	------------------------------------------------------------------------

type machine_state is (

--- generated

ADC_ABSOLUTE_STATE_0,
ADC_ABSOLUTE_STATE_1,
ADC_ABSOLUTE_STATE_2,
ADC_ABSOLUTE_STATE_3,
ADC_ABSOLUTE_STATE_4,
ADC_ABSOLUTE_STATE_5,
ADC_ABSOLUTE_STATE_6,
ADC_ABSOLUTE_STATE_7,
ADC_ABSOLUTE_STATE_8,
ADC_ABSOLUTE_STATE_9,


ADC_ABSOLUTE_X_STATE_0,
ADC_ABSOLUTE_X_STATE_1,
ADC_ABSOLUTE_X_STATE_2,
ADC_ABSOLUTE_X_STATE_3,
ADC_ABSOLUTE_X_STATE_4,
ADC_ABSOLUTE_X_STATE_5,
ADC_ABSOLUTE_X_STATE_6,
ADC_ABSOLUTE_X_STATE_7,
ADC_ABSOLUTE_X_STATE_8,
ADC_ABSOLUTE_X_STATE_9,


ADC_ABSOLUTE_Y_STATE_0,
ADC_ABSOLUTE_Y_STATE_1,
ADC_ABSOLUTE_Y_STATE_2,
ADC_ABSOLUTE_Y_STATE_3,
ADC_ABSOLUTE_Y_STATE_4,
ADC_ABSOLUTE_Y_STATE_5,
ADC_ABSOLUTE_Y_STATE_6,
ADC_ABSOLUTE_Y_STATE_7,
ADC_ABSOLUTE_Y_STATE_8,
ADC_ABSOLUTE_Y_STATE_9,


ADC_IMMEDIATE_STATE_0,
ADC_IMMEDIATE_STATE_1,
ADC_IMMEDIATE_STATE_2,
ADC_IMMEDIATE_STATE_3,
ADC_IMMEDIATE_STATE_4,
ADC_IMMEDIATE_STATE_5,
ADC_IMMEDIATE_STATE_6,
ADC_IMMEDIATE_STATE_7,
ADC_IMMEDIATE_STATE_8,
ADC_IMMEDIATE_STATE_9,


ADC_INDIRECT_X_STATE_0,
ADC_INDIRECT_X_STATE_1,
ADC_INDIRECT_X_STATE_2,
ADC_INDIRECT_X_STATE_3,
ADC_INDIRECT_X_STATE_4,
ADC_INDIRECT_X_STATE_5,
ADC_INDIRECT_X_STATE_6,
ADC_INDIRECT_X_STATE_7,
ADC_INDIRECT_X_STATE_8,
ADC_INDIRECT_X_STATE_9,


ADC_INDIRECT_Y_STATE_0,
ADC_INDIRECT_Y_STATE_1,
ADC_INDIRECT_Y_STATE_2,
ADC_INDIRECT_Y_STATE_3,
ADC_INDIRECT_Y_STATE_4,
ADC_INDIRECT_Y_STATE_5,
ADC_INDIRECT_Y_STATE_6,
ADC_INDIRECT_Y_STATE_7,
ADC_INDIRECT_Y_STATE_8,
ADC_INDIRECT_Y_STATE_9,


ADC_ZERO_PAGE_STATE_0,
ADC_ZERO_PAGE_STATE_1,
ADC_ZERO_PAGE_STATE_2,
ADC_ZERO_PAGE_STATE_3,
ADC_ZERO_PAGE_STATE_4,
ADC_ZERO_PAGE_STATE_5,
ADC_ZERO_PAGE_STATE_6,
ADC_ZERO_PAGE_STATE_7,
ADC_ZERO_PAGE_STATE_8,
ADC_ZERO_PAGE_STATE_9,


ADC_ZERO_PAGE_X_STATE_0,
ADC_ZERO_PAGE_X_STATE_1,
ADC_ZERO_PAGE_X_STATE_2,
ADC_ZERO_PAGE_X_STATE_3,
ADC_ZERO_PAGE_X_STATE_4,
ADC_ZERO_PAGE_X_STATE_5,
ADC_ZERO_PAGE_X_STATE_6,
ADC_ZERO_PAGE_X_STATE_7,
ADC_ZERO_PAGE_X_STATE_8,
ADC_ZERO_PAGE_X_STATE_9,


AND_ABSOLUTE_STATE_0,
AND_ABSOLUTE_STATE_1,
AND_ABSOLUTE_STATE_2,
AND_ABSOLUTE_STATE_3,
AND_ABSOLUTE_STATE_4,
AND_ABSOLUTE_STATE_5,
AND_ABSOLUTE_STATE_6,
AND_ABSOLUTE_STATE_7,
AND_ABSOLUTE_STATE_8,
AND_ABSOLUTE_STATE_9,


AND_ABSOLUTE_X_STATE_0,
AND_ABSOLUTE_X_STATE_1,
AND_ABSOLUTE_X_STATE_2,
AND_ABSOLUTE_X_STATE_3,
AND_ABSOLUTE_X_STATE_4,
AND_ABSOLUTE_X_STATE_5,
AND_ABSOLUTE_X_STATE_6,
AND_ABSOLUTE_X_STATE_7,
AND_ABSOLUTE_X_STATE_8,
AND_ABSOLUTE_X_STATE_9,


AND_ABSOLUTE_Y_STATE_0,
AND_ABSOLUTE_Y_STATE_1,
AND_ABSOLUTE_Y_STATE_2,
AND_ABSOLUTE_Y_STATE_3,
AND_ABSOLUTE_Y_STATE_4,
AND_ABSOLUTE_Y_STATE_5,
AND_ABSOLUTE_Y_STATE_6,
AND_ABSOLUTE_Y_STATE_7,
AND_ABSOLUTE_Y_STATE_8,
AND_ABSOLUTE_Y_STATE_9,


AND_IMMEDIATE_STATE_0,
AND_IMMEDIATE_STATE_1,
AND_IMMEDIATE_STATE_2,
AND_IMMEDIATE_STATE_3,
AND_IMMEDIATE_STATE_4,
AND_IMMEDIATE_STATE_5,
AND_IMMEDIATE_STATE_6,
AND_IMMEDIATE_STATE_7,
AND_IMMEDIATE_STATE_8,
AND_IMMEDIATE_STATE_9,


AND_INDIRECT_X_STATE_0,
AND_INDIRECT_X_STATE_1,
AND_INDIRECT_X_STATE_2,
AND_INDIRECT_X_STATE_3,
AND_INDIRECT_X_STATE_4,
AND_INDIRECT_X_STATE_5,
AND_INDIRECT_X_STATE_6,
AND_INDIRECT_X_STATE_7,
AND_INDIRECT_X_STATE_8,
AND_INDIRECT_X_STATE_9,


AND_INDIRECT_Y_STATE_0,
AND_INDIRECT_Y_STATE_1,
AND_INDIRECT_Y_STATE_2,
AND_INDIRECT_Y_STATE_3,
AND_INDIRECT_Y_STATE_4,
AND_INDIRECT_Y_STATE_5,
AND_INDIRECT_Y_STATE_6,
AND_INDIRECT_Y_STATE_7,
AND_INDIRECT_Y_STATE_8,
AND_INDIRECT_Y_STATE_9,


AND_ZERO_PAGE_STATE_0,
AND_ZERO_PAGE_STATE_1,
AND_ZERO_PAGE_STATE_2,
AND_ZERO_PAGE_STATE_3,
AND_ZERO_PAGE_STATE_4,
AND_ZERO_PAGE_STATE_5,
AND_ZERO_PAGE_STATE_6,
AND_ZERO_PAGE_STATE_7,
AND_ZERO_PAGE_STATE_8,
AND_ZERO_PAGE_STATE_9,


AND_ZERO_PAGE_X_STATE_0,
AND_ZERO_PAGE_X_STATE_1,
AND_ZERO_PAGE_X_STATE_2,
AND_ZERO_PAGE_X_STATE_3,
AND_ZERO_PAGE_X_STATE_4,
AND_ZERO_PAGE_X_STATE_5,
AND_ZERO_PAGE_X_STATE_6,
AND_ZERO_PAGE_X_STATE_7,
AND_ZERO_PAGE_X_STATE_8,
AND_ZERO_PAGE_X_STATE_9,


ASL_ABSOLUTE_STATE_0,
ASL_ABSOLUTE_STATE_1,
ASL_ABSOLUTE_STATE_2,
ASL_ABSOLUTE_STATE_3,
ASL_ABSOLUTE_STATE_4,
ASL_ABSOLUTE_STATE_5,
ASL_ABSOLUTE_STATE_6,
ASL_ABSOLUTE_STATE_7,
ASL_ABSOLUTE_STATE_8,
ASL_ABSOLUTE_STATE_9,


ASL_ABSOLUTE_X_STATE_0,
ASL_ABSOLUTE_X_STATE_1,
ASL_ABSOLUTE_X_STATE_2,
ASL_ABSOLUTE_X_STATE_3,
ASL_ABSOLUTE_X_STATE_4,
ASL_ABSOLUTE_X_STATE_5,
ASL_ABSOLUTE_X_STATE_6,
ASL_ABSOLUTE_X_STATE_7,
ASL_ABSOLUTE_X_STATE_8,
ASL_ABSOLUTE_X_STATE_9,


ASL_ACCUMULATOR_STATE_0,
ASL_ACCUMULATOR_STATE_1,
ASL_ACCUMULATOR_STATE_2,
ASL_ACCUMULATOR_STATE_3,
ASL_ACCUMULATOR_STATE_4,
ASL_ACCUMULATOR_STATE_5,
ASL_ACCUMULATOR_STATE_6,
ASL_ACCUMULATOR_STATE_7,
ASL_ACCUMULATOR_STATE_8,
ASL_ACCUMULATOR_STATE_9,


ASL_ZERO_PAGE_STATE_0,
ASL_ZERO_PAGE_STATE_1,
ASL_ZERO_PAGE_STATE_2,
ASL_ZERO_PAGE_STATE_3,
ASL_ZERO_PAGE_STATE_4,
ASL_ZERO_PAGE_STATE_5,
ASL_ZERO_PAGE_STATE_6,
ASL_ZERO_PAGE_STATE_7,
ASL_ZERO_PAGE_STATE_8,
ASL_ZERO_PAGE_STATE_9,


ASL_ZERO_PAGE_X_STATE_0,
ASL_ZERO_PAGE_X_STATE_1,
ASL_ZERO_PAGE_X_STATE_2,
ASL_ZERO_PAGE_X_STATE_3,
ASL_ZERO_PAGE_X_STATE_4,
ASL_ZERO_PAGE_X_STATE_5,
ASL_ZERO_PAGE_X_STATE_6,
ASL_ZERO_PAGE_X_STATE_7,
ASL_ZERO_PAGE_X_STATE_8,
ASL_ZERO_PAGE_X_STATE_9,


BCC_RELATIVE_STATE_0,
BCC_RELATIVE_STATE_1,
BCC_RELATIVE_STATE_2,
BCC_RELATIVE_STATE_3,
BCC_RELATIVE_STATE_4,
BCC_RELATIVE_STATE_5,
BCC_RELATIVE_STATE_6,
BCC_RELATIVE_STATE_7,
BCC_RELATIVE_STATE_8,
BCC_RELATIVE_STATE_9,


BCS_RELATIVE_STATE_0,
BCS_RELATIVE_STATE_1,
BCS_RELATIVE_STATE_2,
BCS_RELATIVE_STATE_3,
BCS_RELATIVE_STATE_4,
BCS_RELATIVE_STATE_5,
BCS_RELATIVE_STATE_6,
BCS_RELATIVE_STATE_7,
BCS_RELATIVE_STATE_8,
BCS_RELATIVE_STATE_9,


BEQ_RELATIVE_STATE_0,
BEQ_RELATIVE_STATE_1,
BEQ_RELATIVE_STATE_2,
BEQ_RELATIVE_STATE_3,
BEQ_RELATIVE_STATE_4,
BEQ_RELATIVE_STATE_5,
BEQ_RELATIVE_STATE_6,
BEQ_RELATIVE_STATE_7,
BEQ_RELATIVE_STATE_8,
BEQ_RELATIVE_STATE_9,


BIT_ABSOLUTE_STATE_0,
BIT_ABSOLUTE_STATE_1,
BIT_ABSOLUTE_STATE_2,
BIT_ABSOLUTE_STATE_3,
BIT_ABSOLUTE_STATE_4,
BIT_ABSOLUTE_STATE_5,
BIT_ABSOLUTE_STATE_6,
BIT_ABSOLUTE_STATE_7,
BIT_ABSOLUTE_STATE_8,
BIT_ABSOLUTE_STATE_9,


BIT_ZERO_PAGE_STATE_0,
BIT_ZERO_PAGE_STATE_1,
BIT_ZERO_PAGE_STATE_2,
BIT_ZERO_PAGE_STATE_3,
BIT_ZERO_PAGE_STATE_4,
BIT_ZERO_PAGE_STATE_5,
BIT_ZERO_PAGE_STATE_6,
BIT_ZERO_PAGE_STATE_7,
BIT_ZERO_PAGE_STATE_8,
BIT_ZERO_PAGE_STATE_9,


BMI_RELATIVE_STATE_0,
BMI_RELATIVE_STATE_1,
BMI_RELATIVE_STATE_2,
BMI_RELATIVE_STATE_3,
BMI_RELATIVE_STATE_4,
BMI_RELATIVE_STATE_5,
BMI_RELATIVE_STATE_6,
BMI_RELATIVE_STATE_7,
BMI_RELATIVE_STATE_8,
BMI_RELATIVE_STATE_9,


BNE_RELATIVE_STATE_0,
BNE_RELATIVE_STATE_1,
BNE_RELATIVE_STATE_2,
BNE_RELATIVE_STATE_3,
BNE_RELATIVE_STATE_4,
BNE_RELATIVE_STATE_5,
BNE_RELATIVE_STATE_6,
BNE_RELATIVE_STATE_7,
BNE_RELATIVE_STATE_8,
BNE_RELATIVE_STATE_9,


BPL_RELATIVE_STATE_0,
BPL_RELATIVE_STATE_1,
BPL_RELATIVE_STATE_2,
BPL_RELATIVE_STATE_3,
BPL_RELATIVE_STATE_4,
BPL_RELATIVE_STATE_5,
BPL_RELATIVE_STATE_6,
BPL_RELATIVE_STATE_7,
BPL_RELATIVE_STATE_8,
BPL_RELATIVE_STATE_9,


BRK_IMPLIED_STATE_0,
BRK_IMPLIED_STATE_1,
BRK_IMPLIED_STATE_2,
BRK_IMPLIED_STATE_3,
BRK_IMPLIED_STATE_4,
BRK_IMPLIED_STATE_5,
BRK_IMPLIED_STATE_6,
BRK_IMPLIED_STATE_7,
BRK_IMPLIED_STATE_8,
BRK_IMPLIED_STATE_9,


BVC_RELATIVE_STATE_0,
BVC_RELATIVE_STATE_1,
BVC_RELATIVE_STATE_2,
BVC_RELATIVE_STATE_3,
BVC_RELATIVE_STATE_4,
BVC_RELATIVE_STATE_5,
BVC_RELATIVE_STATE_6,
BVC_RELATIVE_STATE_7,
BVC_RELATIVE_STATE_8,
BVC_RELATIVE_STATE_9,


BVS_RELATIVE_STATE_0,
BVS_RELATIVE_STATE_1,
BVS_RELATIVE_STATE_2,
BVS_RELATIVE_STATE_3,
BVS_RELATIVE_STATE_4,
BVS_RELATIVE_STATE_5,
BVS_RELATIVE_STATE_6,
BVS_RELATIVE_STATE_7,
BVS_RELATIVE_STATE_8,
BVS_RELATIVE_STATE_9,


CLC_IMPLIED_STATE_0,
CLC_IMPLIED_STATE_1,
CLC_IMPLIED_STATE_2,
CLC_IMPLIED_STATE_3,
CLC_IMPLIED_STATE_4,
CLC_IMPLIED_STATE_5,
CLC_IMPLIED_STATE_6,
CLC_IMPLIED_STATE_7,
CLC_IMPLIED_STATE_8,
CLC_IMPLIED_STATE_9,


CLD_IMPLIED_STATE_0,
CLD_IMPLIED_STATE_1,
CLD_IMPLIED_STATE_2,
CLD_IMPLIED_STATE_3,
CLD_IMPLIED_STATE_4,
CLD_IMPLIED_STATE_5,
CLD_IMPLIED_STATE_6,
CLD_IMPLIED_STATE_7,
CLD_IMPLIED_STATE_8,
CLD_IMPLIED_STATE_9,


CLI_IMPLIED_STATE_0,
CLI_IMPLIED_STATE_1,
CLI_IMPLIED_STATE_2,
CLI_IMPLIED_STATE_3,
CLI_IMPLIED_STATE_4,
CLI_IMPLIED_STATE_5,
CLI_IMPLIED_STATE_6,
CLI_IMPLIED_STATE_7,
CLI_IMPLIED_STATE_8,
CLI_IMPLIED_STATE_9,


CLV_IMPLIED_STATE_0,
CLV_IMPLIED_STATE_1,
CLV_IMPLIED_STATE_2,
CLV_IMPLIED_STATE_3,
CLV_IMPLIED_STATE_4,
CLV_IMPLIED_STATE_5,
CLV_IMPLIED_STATE_6,
CLV_IMPLIED_STATE_7,
CLV_IMPLIED_STATE_8,
CLV_IMPLIED_STATE_9,


CMP_ABSOLUTE_STATE_0,
CMP_ABSOLUTE_STATE_1,
CMP_ABSOLUTE_STATE_2,
CMP_ABSOLUTE_STATE_3,
CMP_ABSOLUTE_STATE_4,
CMP_ABSOLUTE_STATE_5,
CMP_ABSOLUTE_STATE_6,
CMP_ABSOLUTE_STATE_7,
CMP_ABSOLUTE_STATE_8,
CMP_ABSOLUTE_STATE_9,


CMP_ABSOLUTE_X_STATE_0,
CMP_ABSOLUTE_X_STATE_1,
CMP_ABSOLUTE_X_STATE_2,
CMP_ABSOLUTE_X_STATE_3,
CMP_ABSOLUTE_X_STATE_4,
CMP_ABSOLUTE_X_STATE_5,
CMP_ABSOLUTE_X_STATE_6,
CMP_ABSOLUTE_X_STATE_7,
CMP_ABSOLUTE_X_STATE_8,
CMP_ABSOLUTE_X_STATE_9,


CMP_ABSOLUTE_Y_STATE_0,
CMP_ABSOLUTE_Y_STATE_1,
CMP_ABSOLUTE_Y_STATE_2,
CMP_ABSOLUTE_Y_STATE_3,
CMP_ABSOLUTE_Y_STATE_4,
CMP_ABSOLUTE_Y_STATE_5,
CMP_ABSOLUTE_Y_STATE_6,
CMP_ABSOLUTE_Y_STATE_7,
CMP_ABSOLUTE_Y_STATE_8,
CMP_ABSOLUTE_Y_STATE_9,


CMP_IMMEDIATE_STATE_0,
CMP_IMMEDIATE_STATE_1,
CMP_IMMEDIATE_STATE_2,
CMP_IMMEDIATE_STATE_3,
CMP_IMMEDIATE_STATE_4,
CMP_IMMEDIATE_STATE_5,
CMP_IMMEDIATE_STATE_6,
CMP_IMMEDIATE_STATE_7,
CMP_IMMEDIATE_STATE_8,
CMP_IMMEDIATE_STATE_9,


CMP_INDIRECT_X_STATE_0,
CMP_INDIRECT_X_STATE_1,
CMP_INDIRECT_X_STATE_2,
CMP_INDIRECT_X_STATE_3,
CMP_INDIRECT_X_STATE_4,
CMP_INDIRECT_X_STATE_5,
CMP_INDIRECT_X_STATE_6,
CMP_INDIRECT_X_STATE_7,
CMP_INDIRECT_X_STATE_8,
CMP_INDIRECT_X_STATE_9,


CMP_INDIRECT_Y_STATE_0,
CMP_INDIRECT_Y_STATE_1,
CMP_INDIRECT_Y_STATE_2,
CMP_INDIRECT_Y_STATE_3,
CMP_INDIRECT_Y_STATE_4,
CMP_INDIRECT_Y_STATE_5,
CMP_INDIRECT_Y_STATE_6,
CMP_INDIRECT_Y_STATE_7,
CMP_INDIRECT_Y_STATE_8,
CMP_INDIRECT_Y_STATE_9,


CMP_ZERO_PAGE_STATE_0,
CMP_ZERO_PAGE_STATE_1,
CMP_ZERO_PAGE_STATE_2,
CMP_ZERO_PAGE_STATE_3,
CMP_ZERO_PAGE_STATE_4,
CMP_ZERO_PAGE_STATE_5,
CMP_ZERO_PAGE_STATE_6,
CMP_ZERO_PAGE_STATE_7,
CMP_ZERO_PAGE_STATE_8,
CMP_ZERO_PAGE_STATE_9,


CMP_ZERO_PAGE_X_STATE_0,
CMP_ZERO_PAGE_X_STATE_1,
CMP_ZERO_PAGE_X_STATE_2,
CMP_ZERO_PAGE_X_STATE_3,
CMP_ZERO_PAGE_X_STATE_4,
CMP_ZERO_PAGE_X_STATE_5,
CMP_ZERO_PAGE_X_STATE_6,
CMP_ZERO_PAGE_X_STATE_7,
CMP_ZERO_PAGE_X_STATE_8,
CMP_ZERO_PAGE_X_STATE_9,


CPX_ABSOLUTE_STATE_0,
CPX_ABSOLUTE_STATE_1,
CPX_ABSOLUTE_STATE_2,
CPX_ABSOLUTE_STATE_3,
CPX_ABSOLUTE_STATE_4,
CPX_ABSOLUTE_STATE_5,
CPX_ABSOLUTE_STATE_6,
CPX_ABSOLUTE_STATE_7,
CPX_ABSOLUTE_STATE_8,
CPX_ABSOLUTE_STATE_9,


CPX_IMMEDIATE_STATE_0,
CPX_IMMEDIATE_STATE_1,
CPX_IMMEDIATE_STATE_2,
CPX_IMMEDIATE_STATE_3,
CPX_IMMEDIATE_STATE_4,
CPX_IMMEDIATE_STATE_5,
CPX_IMMEDIATE_STATE_6,
CPX_IMMEDIATE_STATE_7,
CPX_IMMEDIATE_STATE_8,
CPX_IMMEDIATE_STATE_9,


CPX_ZERO_PAGE_STATE_0,
CPX_ZERO_PAGE_STATE_1,
CPX_ZERO_PAGE_STATE_2,
CPX_ZERO_PAGE_STATE_3,
CPX_ZERO_PAGE_STATE_4,
CPX_ZERO_PAGE_STATE_5,
CPX_ZERO_PAGE_STATE_6,
CPX_ZERO_PAGE_STATE_7,
CPX_ZERO_PAGE_STATE_8,
CPX_ZERO_PAGE_STATE_9,


CPY_ABSOLUTE_STATE_0,
CPY_ABSOLUTE_STATE_1,
CPY_ABSOLUTE_STATE_2,
CPY_ABSOLUTE_STATE_3,
CPY_ABSOLUTE_STATE_4,
CPY_ABSOLUTE_STATE_5,
CPY_ABSOLUTE_STATE_6,
CPY_ABSOLUTE_STATE_7,
CPY_ABSOLUTE_STATE_8,
CPY_ABSOLUTE_STATE_9,


CPY_IMMEDIATE_STATE_0,
CPY_IMMEDIATE_STATE_1,
CPY_IMMEDIATE_STATE_2,
CPY_IMMEDIATE_STATE_3,
CPY_IMMEDIATE_STATE_4,
CPY_IMMEDIATE_STATE_5,
CPY_IMMEDIATE_STATE_6,
CPY_IMMEDIATE_STATE_7,
CPY_IMMEDIATE_STATE_8,
CPY_IMMEDIATE_STATE_9,


CPY_ZERO_PAGE_STATE_0,
CPY_ZERO_PAGE_STATE_1,
CPY_ZERO_PAGE_STATE_2,
CPY_ZERO_PAGE_STATE_3,
CPY_ZERO_PAGE_STATE_4,
CPY_ZERO_PAGE_STATE_5,
CPY_ZERO_PAGE_STATE_6,
CPY_ZERO_PAGE_STATE_7,
CPY_ZERO_PAGE_STATE_8,
CPY_ZERO_PAGE_STATE_9,


DEC_ABSOLUTE_STATE_0,
DEC_ABSOLUTE_STATE_1,
DEC_ABSOLUTE_STATE_2,
DEC_ABSOLUTE_STATE_3,
DEC_ABSOLUTE_STATE_4,
DEC_ABSOLUTE_STATE_5,
DEC_ABSOLUTE_STATE_6,
DEC_ABSOLUTE_STATE_7,
DEC_ABSOLUTE_STATE_8,
DEC_ABSOLUTE_STATE_9,


DEC_ABSOLUTE_X_STATE_0,
DEC_ABSOLUTE_X_STATE_1,
DEC_ABSOLUTE_X_STATE_2,
DEC_ABSOLUTE_X_STATE_3,
DEC_ABSOLUTE_X_STATE_4,
DEC_ABSOLUTE_X_STATE_5,
DEC_ABSOLUTE_X_STATE_6,
DEC_ABSOLUTE_X_STATE_7,
DEC_ABSOLUTE_X_STATE_8,
DEC_ABSOLUTE_X_STATE_9,


DEC_ZERO_PAGE_STATE_0,
DEC_ZERO_PAGE_STATE_1,
DEC_ZERO_PAGE_STATE_2,
DEC_ZERO_PAGE_STATE_3,
DEC_ZERO_PAGE_STATE_4,
DEC_ZERO_PAGE_STATE_5,
DEC_ZERO_PAGE_STATE_6,
DEC_ZERO_PAGE_STATE_7,
DEC_ZERO_PAGE_STATE_8,
DEC_ZERO_PAGE_STATE_9,


DEC_ZERO_PAGE_X_STATE_0,
DEC_ZERO_PAGE_X_STATE_1,
DEC_ZERO_PAGE_X_STATE_2,
DEC_ZERO_PAGE_X_STATE_3,
DEC_ZERO_PAGE_X_STATE_4,
DEC_ZERO_PAGE_X_STATE_5,
DEC_ZERO_PAGE_X_STATE_6,
DEC_ZERO_PAGE_X_STATE_7,
DEC_ZERO_PAGE_X_STATE_8,
DEC_ZERO_PAGE_X_STATE_9,


DEX_IMPLIED_STATE_0,
DEX_IMPLIED_STATE_1,
DEX_IMPLIED_STATE_2,
DEX_IMPLIED_STATE_3,
DEX_IMPLIED_STATE_4,
DEX_IMPLIED_STATE_5,
DEX_IMPLIED_STATE_6,
DEX_IMPLIED_STATE_7,
DEX_IMPLIED_STATE_8,
DEX_IMPLIED_STATE_9,


DEY_IMPLIED_STATE_0,
DEY_IMPLIED_STATE_1,
DEY_IMPLIED_STATE_2,
DEY_IMPLIED_STATE_3,
DEY_IMPLIED_STATE_4,
DEY_IMPLIED_STATE_5,
DEY_IMPLIED_STATE_6,
DEY_IMPLIED_STATE_7,
DEY_IMPLIED_STATE_8,
DEY_IMPLIED_STATE_9,


EOR_ABSOLUTE_STATE_0,
EOR_ABSOLUTE_STATE_1,
EOR_ABSOLUTE_STATE_2,
EOR_ABSOLUTE_STATE_3,
EOR_ABSOLUTE_STATE_4,
EOR_ABSOLUTE_STATE_5,
EOR_ABSOLUTE_STATE_6,
EOR_ABSOLUTE_STATE_7,
EOR_ABSOLUTE_STATE_8,
EOR_ABSOLUTE_STATE_9,


EOR_ABSOLUTE_X_STATE_0,
EOR_ABSOLUTE_X_STATE_1,
EOR_ABSOLUTE_X_STATE_2,
EOR_ABSOLUTE_X_STATE_3,
EOR_ABSOLUTE_X_STATE_4,
EOR_ABSOLUTE_X_STATE_5,
EOR_ABSOLUTE_X_STATE_6,
EOR_ABSOLUTE_X_STATE_7,
EOR_ABSOLUTE_X_STATE_8,
EOR_ABSOLUTE_X_STATE_9,


EOR_ABSOLUTE_Y_STATE_0,
EOR_ABSOLUTE_Y_STATE_1,
EOR_ABSOLUTE_Y_STATE_2,
EOR_ABSOLUTE_Y_STATE_3,
EOR_ABSOLUTE_Y_STATE_4,
EOR_ABSOLUTE_Y_STATE_5,
EOR_ABSOLUTE_Y_STATE_6,
EOR_ABSOLUTE_Y_STATE_7,
EOR_ABSOLUTE_Y_STATE_8,
EOR_ABSOLUTE_Y_STATE_9,


EOR_IMMEDIATE_STATE_0,
EOR_IMMEDIATE_STATE_1,
EOR_IMMEDIATE_STATE_2,
EOR_IMMEDIATE_STATE_3,
EOR_IMMEDIATE_STATE_4,
EOR_IMMEDIATE_STATE_5,
EOR_IMMEDIATE_STATE_6,
EOR_IMMEDIATE_STATE_7,
EOR_IMMEDIATE_STATE_8,
EOR_IMMEDIATE_STATE_9,


EOR_INDIRECT_X_STATE_0,
EOR_INDIRECT_X_STATE_1,
EOR_INDIRECT_X_STATE_2,
EOR_INDIRECT_X_STATE_3,
EOR_INDIRECT_X_STATE_4,
EOR_INDIRECT_X_STATE_5,
EOR_INDIRECT_X_STATE_6,
EOR_INDIRECT_X_STATE_7,
EOR_INDIRECT_X_STATE_8,
EOR_INDIRECT_X_STATE_9,


EOR_INDIRECT_Y_STATE_0,
EOR_INDIRECT_Y_STATE_1,
EOR_INDIRECT_Y_STATE_2,
EOR_INDIRECT_Y_STATE_3,
EOR_INDIRECT_Y_STATE_4,
EOR_INDIRECT_Y_STATE_5,
EOR_INDIRECT_Y_STATE_6,
EOR_INDIRECT_Y_STATE_7,
EOR_INDIRECT_Y_STATE_8,
EOR_INDIRECT_Y_STATE_9,


EOR_ZERO_PAGE_STATE_0,
EOR_ZERO_PAGE_STATE_1,
EOR_ZERO_PAGE_STATE_2,
EOR_ZERO_PAGE_STATE_3,
EOR_ZERO_PAGE_STATE_4,
EOR_ZERO_PAGE_STATE_5,
EOR_ZERO_PAGE_STATE_6,
EOR_ZERO_PAGE_STATE_7,
EOR_ZERO_PAGE_STATE_8,
EOR_ZERO_PAGE_STATE_9,


EOR_ZERO_PAGE_X_STATE_0,
EOR_ZERO_PAGE_X_STATE_1,
EOR_ZERO_PAGE_X_STATE_2,
EOR_ZERO_PAGE_X_STATE_3,
EOR_ZERO_PAGE_X_STATE_4,
EOR_ZERO_PAGE_X_STATE_5,
EOR_ZERO_PAGE_X_STATE_6,
EOR_ZERO_PAGE_X_STATE_7,
EOR_ZERO_PAGE_X_STATE_8,
EOR_ZERO_PAGE_X_STATE_9,


INC_ABSOLUTE_STATE_0,
INC_ABSOLUTE_STATE_1,
INC_ABSOLUTE_STATE_2,
INC_ABSOLUTE_STATE_3,
INC_ABSOLUTE_STATE_4,
INC_ABSOLUTE_STATE_5,
INC_ABSOLUTE_STATE_6,
INC_ABSOLUTE_STATE_7,
INC_ABSOLUTE_STATE_8,
INC_ABSOLUTE_STATE_9,


INC_ABSOLUTE_X_STATE_0,
INC_ABSOLUTE_X_STATE_1,
INC_ABSOLUTE_X_STATE_2,
INC_ABSOLUTE_X_STATE_3,
INC_ABSOLUTE_X_STATE_4,
INC_ABSOLUTE_X_STATE_5,
INC_ABSOLUTE_X_STATE_6,
INC_ABSOLUTE_X_STATE_7,
INC_ABSOLUTE_X_STATE_8,
INC_ABSOLUTE_X_STATE_9,


INC_ZERO_PAGE_STATE_0,
INC_ZERO_PAGE_STATE_1,
INC_ZERO_PAGE_STATE_2,
INC_ZERO_PAGE_STATE_3,
INC_ZERO_PAGE_STATE_4,
INC_ZERO_PAGE_STATE_5,
INC_ZERO_PAGE_STATE_6,
INC_ZERO_PAGE_STATE_7,
INC_ZERO_PAGE_STATE_8,
INC_ZERO_PAGE_STATE_9,


INC_ZERO_PAGE_X_STATE_0,
INC_ZERO_PAGE_X_STATE_1,
INC_ZERO_PAGE_X_STATE_2,
INC_ZERO_PAGE_X_STATE_3,
INC_ZERO_PAGE_X_STATE_4,
INC_ZERO_PAGE_X_STATE_5,
INC_ZERO_PAGE_X_STATE_6,
INC_ZERO_PAGE_X_STATE_7,
INC_ZERO_PAGE_X_STATE_8,
INC_ZERO_PAGE_X_STATE_9,


INX_IMPLIED_STATE_0,
INX_IMPLIED_STATE_1,
INX_IMPLIED_STATE_2,
INX_IMPLIED_STATE_3,
INX_IMPLIED_STATE_4,
INX_IMPLIED_STATE_5,
INX_IMPLIED_STATE_6,
INX_IMPLIED_STATE_7,
INX_IMPLIED_STATE_8,
INX_IMPLIED_STATE_9,


INY_IMPLIED_STATE_0,
INY_IMPLIED_STATE_1,
INY_IMPLIED_STATE_2,
INY_IMPLIED_STATE_3,
INY_IMPLIED_STATE_4,
INY_IMPLIED_STATE_5,
INY_IMPLIED_STATE_6,
INY_IMPLIED_STATE_7,
INY_IMPLIED_STATE_8,
INY_IMPLIED_STATE_9,


JMP_ABSOLUTE_STATE_0,
JMP_ABSOLUTE_STATE_1,
JMP_ABSOLUTE_STATE_2,
JMP_ABSOLUTE_STATE_3,
JMP_ABSOLUTE_STATE_4,
JMP_ABSOLUTE_STATE_5,
JMP_ABSOLUTE_STATE_6,
JMP_ABSOLUTE_STATE_7,
JMP_ABSOLUTE_STATE_8,
JMP_ABSOLUTE_STATE_9,


JMP_INDIRECT_STATE_0,
JMP_INDIRECT_STATE_1,
JMP_INDIRECT_STATE_2,
JMP_INDIRECT_STATE_3,
JMP_INDIRECT_STATE_4,
JMP_INDIRECT_STATE_5,
JMP_INDIRECT_STATE_6,
JMP_INDIRECT_STATE_7,
JMP_INDIRECT_STATE_8,
JMP_INDIRECT_STATE_9,


JSR_ABSOLUTE_STATE_0,
JSR_ABSOLUTE_STATE_1,
JSR_ABSOLUTE_STATE_2,
JSR_ABSOLUTE_STATE_3,
JSR_ABSOLUTE_STATE_4,
JSR_ABSOLUTE_STATE_5,
JSR_ABSOLUTE_STATE_6,
JSR_ABSOLUTE_STATE_7,
JSR_ABSOLUTE_STATE_8,
JSR_ABSOLUTE_STATE_9,


LDA_ABSOLUTE_STATE_0,
LDA_ABSOLUTE_STATE_1,
LDA_ABSOLUTE_STATE_2,
LDA_ABSOLUTE_STATE_3,
LDA_ABSOLUTE_STATE_4,
LDA_ABSOLUTE_STATE_5,
LDA_ABSOLUTE_STATE_6,
LDA_ABSOLUTE_STATE_7,
LDA_ABSOLUTE_STATE_8,
LDA_ABSOLUTE_STATE_9,


LDA_ABSOLUTE_X_STATE_0,
LDA_ABSOLUTE_X_STATE_1,
LDA_ABSOLUTE_X_STATE_2,
LDA_ABSOLUTE_X_STATE_3,
LDA_ABSOLUTE_X_STATE_4,
LDA_ABSOLUTE_X_STATE_5,
LDA_ABSOLUTE_X_STATE_6,
LDA_ABSOLUTE_X_STATE_7,
LDA_ABSOLUTE_X_STATE_8,
LDA_ABSOLUTE_X_STATE_9,


LDA_ABSOLUTE_Y_STATE_0,
LDA_ABSOLUTE_Y_STATE_1,
LDA_ABSOLUTE_Y_STATE_2,
LDA_ABSOLUTE_Y_STATE_3,
LDA_ABSOLUTE_Y_STATE_4,
LDA_ABSOLUTE_Y_STATE_5,
LDA_ABSOLUTE_Y_STATE_6,
LDA_ABSOLUTE_Y_STATE_7,
LDA_ABSOLUTE_Y_STATE_8,
LDA_ABSOLUTE_Y_STATE_9,


LDA_IMMEDIATE_STATE_0,
LDA_IMMEDIATE_STATE_1,
LDA_IMMEDIATE_STATE_2,
LDA_IMMEDIATE_STATE_3,
LDA_IMMEDIATE_STATE_4,
LDA_IMMEDIATE_STATE_5,
LDA_IMMEDIATE_STATE_6,
LDA_IMMEDIATE_STATE_7,
LDA_IMMEDIATE_STATE_8,
LDA_IMMEDIATE_STATE_9,


LDA_ZERO_PAGE_STATE_0,
LDA_ZERO_PAGE_STATE_1,
LDA_ZERO_PAGE_STATE_2,
LDA_ZERO_PAGE_STATE_3,
LDA_ZERO_PAGE_STATE_4,
LDA_ZERO_PAGE_STATE_5,
LDA_ZERO_PAGE_STATE_6,
LDA_ZERO_PAGE_STATE_7,
LDA_ZERO_PAGE_STATE_8,
LDA_ZERO_PAGE_STATE_9,


LDA_INDIRECT_X_STATE_0,
LDA_INDIRECT_X_STATE_1,
LDA_INDIRECT_X_STATE_2,
LDA_INDIRECT_X_STATE_3,
LDA_INDIRECT_X_STATE_4,
LDA_INDIRECT_X_STATE_5,
LDA_INDIRECT_X_STATE_6,
LDA_INDIRECT_X_STATE_7,
LDA_INDIRECT_X_STATE_8,
LDA_INDIRECT_X_STATE_9,


LDA_INDIRECT_Y_STATE_0,
LDA_INDIRECT_Y_STATE_1,
LDA_INDIRECT_Y_STATE_2,
LDA_INDIRECT_Y_STATE_3,
LDA_INDIRECT_Y_STATE_4,
LDA_INDIRECT_Y_STATE_5,
LDA_INDIRECT_Y_STATE_6,
LDA_INDIRECT_Y_STATE_7,
LDA_INDIRECT_Y_STATE_8,
LDA_INDIRECT_Y_STATE_9,


LDA_ZERO_PAGE_X_STATE_0,
LDA_ZERO_PAGE_X_STATE_1,
LDA_ZERO_PAGE_X_STATE_2,
LDA_ZERO_PAGE_X_STATE_3,
LDA_ZERO_PAGE_X_STATE_4,
LDA_ZERO_PAGE_X_STATE_5,
LDA_ZERO_PAGE_X_STATE_6,
LDA_ZERO_PAGE_X_STATE_7,
LDA_ZERO_PAGE_X_STATE_8,
LDA_ZERO_PAGE_X_STATE_9,


LDX_ABSOLUTE_STATE_0,
LDX_ABSOLUTE_STATE_1,
LDX_ABSOLUTE_STATE_2,
LDX_ABSOLUTE_STATE_3,
LDX_ABSOLUTE_STATE_4,
LDX_ABSOLUTE_STATE_5,
LDX_ABSOLUTE_STATE_6,
LDX_ABSOLUTE_STATE_7,
LDX_ABSOLUTE_STATE_8,
LDX_ABSOLUTE_STATE_9,


LDX_ABSOLUTE_Y_STATE_0,
LDX_ABSOLUTE_Y_STATE_1,
LDX_ABSOLUTE_Y_STATE_2,
LDX_ABSOLUTE_Y_STATE_3,
LDX_ABSOLUTE_Y_STATE_4,
LDX_ABSOLUTE_Y_STATE_5,
LDX_ABSOLUTE_Y_STATE_6,
LDX_ABSOLUTE_Y_STATE_7,
LDX_ABSOLUTE_Y_STATE_8,
LDX_ABSOLUTE_Y_STATE_9,


LDX_IMMEDIATE_STATE_0,
LDX_IMMEDIATE_STATE_1,
LDX_IMMEDIATE_STATE_2,
LDX_IMMEDIATE_STATE_3,
LDX_IMMEDIATE_STATE_4,
LDX_IMMEDIATE_STATE_5,
LDX_IMMEDIATE_STATE_6,
LDX_IMMEDIATE_STATE_7,
LDX_IMMEDIATE_STATE_8,
LDX_IMMEDIATE_STATE_9,


LDX_ZERO_PAGE_STATE_0,
LDX_ZERO_PAGE_STATE_1,
LDX_ZERO_PAGE_STATE_2,
LDX_ZERO_PAGE_STATE_3,
LDX_ZERO_PAGE_STATE_4,
LDX_ZERO_PAGE_STATE_5,
LDX_ZERO_PAGE_STATE_6,
LDX_ZERO_PAGE_STATE_7,
LDX_ZERO_PAGE_STATE_8,
LDX_ZERO_PAGE_STATE_9,


LDX_ZERO_PAGE_Y_STATE_0,
LDX_ZERO_PAGE_Y_STATE_1,
LDX_ZERO_PAGE_Y_STATE_2,
LDX_ZERO_PAGE_Y_STATE_3,
LDX_ZERO_PAGE_Y_STATE_4,
LDX_ZERO_PAGE_Y_STATE_5,
LDX_ZERO_PAGE_Y_STATE_6,
LDX_ZERO_PAGE_Y_STATE_7,
LDX_ZERO_PAGE_Y_STATE_8,
LDX_ZERO_PAGE_Y_STATE_9,


LDY_ABSOLUTE_STATE_0,
LDY_ABSOLUTE_STATE_1,
LDY_ABSOLUTE_STATE_2,
LDY_ABSOLUTE_STATE_3,
LDY_ABSOLUTE_STATE_4,
LDY_ABSOLUTE_STATE_5,
LDY_ABSOLUTE_STATE_6,
LDY_ABSOLUTE_STATE_7,
LDY_ABSOLUTE_STATE_8,
LDY_ABSOLUTE_STATE_9,


LDY_ABSOLUTE_X_STATE_0,
LDY_ABSOLUTE_X_STATE_1,
LDY_ABSOLUTE_X_STATE_2,
LDY_ABSOLUTE_X_STATE_3,
LDY_ABSOLUTE_X_STATE_4,
LDY_ABSOLUTE_X_STATE_5,
LDY_ABSOLUTE_X_STATE_6,
LDY_ABSOLUTE_X_STATE_7,
LDY_ABSOLUTE_X_STATE_8,
LDY_ABSOLUTE_X_STATE_9,


LDY_IMMEDIATE_STATE_0,
LDY_IMMEDIATE_STATE_1,
LDY_IMMEDIATE_STATE_2,
LDY_IMMEDIATE_STATE_3,
LDY_IMMEDIATE_STATE_4,
LDY_IMMEDIATE_STATE_5,
LDY_IMMEDIATE_STATE_6,
LDY_IMMEDIATE_STATE_7,
LDY_IMMEDIATE_STATE_8,
LDY_IMMEDIATE_STATE_9,


LDY_ZERO_PAGE_STATE_0,
LDY_ZERO_PAGE_STATE_1,
LDY_ZERO_PAGE_STATE_2,
LDY_ZERO_PAGE_STATE_3,
LDY_ZERO_PAGE_STATE_4,
LDY_ZERO_PAGE_STATE_5,
LDY_ZERO_PAGE_STATE_6,
LDY_ZERO_PAGE_STATE_7,
LDY_ZERO_PAGE_STATE_8,
LDY_ZERO_PAGE_STATE_9,


LDY_ZERO_PAGE_X_STATE_0,
LDY_ZERO_PAGE_X_STATE_1,
LDY_ZERO_PAGE_X_STATE_2,
LDY_ZERO_PAGE_X_STATE_3,
LDY_ZERO_PAGE_X_STATE_4,
LDY_ZERO_PAGE_X_STATE_5,
LDY_ZERO_PAGE_X_STATE_6,
LDY_ZERO_PAGE_X_STATE_7,
LDY_ZERO_PAGE_X_STATE_8,
LDY_ZERO_PAGE_X_STATE_9,


LSR_ABSOLUTE_STATE_0,
LSR_ABSOLUTE_STATE_1,
LSR_ABSOLUTE_STATE_2,
LSR_ABSOLUTE_STATE_3,
LSR_ABSOLUTE_STATE_4,
LSR_ABSOLUTE_STATE_5,
LSR_ABSOLUTE_STATE_6,
LSR_ABSOLUTE_STATE_7,
LSR_ABSOLUTE_STATE_8,
LSR_ABSOLUTE_STATE_9,


LSR_ABSOLUTE_X_STATE_0,
LSR_ABSOLUTE_X_STATE_1,
LSR_ABSOLUTE_X_STATE_2,
LSR_ABSOLUTE_X_STATE_3,
LSR_ABSOLUTE_X_STATE_4,
LSR_ABSOLUTE_X_STATE_5,
LSR_ABSOLUTE_X_STATE_6,
LSR_ABSOLUTE_X_STATE_7,
LSR_ABSOLUTE_X_STATE_8,
LSR_ABSOLUTE_X_STATE_9,


LSR_ACCUMULATOR_STATE_0,
LSR_ACCUMULATOR_STATE_1,
LSR_ACCUMULATOR_STATE_2,
LSR_ACCUMULATOR_STATE_3,
LSR_ACCUMULATOR_STATE_4,
LSR_ACCUMULATOR_STATE_5,
LSR_ACCUMULATOR_STATE_6,
LSR_ACCUMULATOR_STATE_7,
LSR_ACCUMULATOR_STATE_8,
LSR_ACCUMULATOR_STATE_9,


LSR_ZERO_PAGE_STATE_0,
LSR_ZERO_PAGE_STATE_1,
LSR_ZERO_PAGE_STATE_2,
LSR_ZERO_PAGE_STATE_3,
LSR_ZERO_PAGE_STATE_4,
LSR_ZERO_PAGE_STATE_5,
LSR_ZERO_PAGE_STATE_6,
LSR_ZERO_PAGE_STATE_7,
LSR_ZERO_PAGE_STATE_8,
LSR_ZERO_PAGE_STATE_9,


LSR_ZERO_PAGE_X_STATE_0,
LSR_ZERO_PAGE_X_STATE_1,
LSR_ZERO_PAGE_X_STATE_2,
LSR_ZERO_PAGE_X_STATE_3,
LSR_ZERO_PAGE_X_STATE_4,
LSR_ZERO_PAGE_X_STATE_5,
LSR_ZERO_PAGE_X_STATE_6,
LSR_ZERO_PAGE_X_STATE_7,
LSR_ZERO_PAGE_X_STATE_8,
LSR_ZERO_PAGE_X_STATE_9,


NOP_IMPLIED_STATE_0,
NOP_IMPLIED_STATE_1,
NOP_IMPLIED_STATE_2,
NOP_IMPLIED_STATE_3,
NOP_IMPLIED_STATE_4,
NOP_IMPLIED_STATE_5,
NOP_IMPLIED_STATE_6,
NOP_IMPLIED_STATE_7,
NOP_IMPLIED_STATE_8,
NOP_IMPLIED_STATE_9,


ORA_ABSOLUTE_STATE_0,
ORA_ABSOLUTE_STATE_1,
ORA_ABSOLUTE_STATE_2,
ORA_ABSOLUTE_STATE_3,
ORA_ABSOLUTE_STATE_4,
ORA_ABSOLUTE_STATE_5,
ORA_ABSOLUTE_STATE_6,
ORA_ABSOLUTE_STATE_7,
ORA_ABSOLUTE_STATE_8,
ORA_ABSOLUTE_STATE_9,


ORA_ABSOLUTE_X_STATE_0,
ORA_ABSOLUTE_X_STATE_1,
ORA_ABSOLUTE_X_STATE_2,
ORA_ABSOLUTE_X_STATE_3,
ORA_ABSOLUTE_X_STATE_4,
ORA_ABSOLUTE_X_STATE_5,
ORA_ABSOLUTE_X_STATE_6,
ORA_ABSOLUTE_X_STATE_7,
ORA_ABSOLUTE_X_STATE_8,
ORA_ABSOLUTE_X_STATE_9,


ORA_ABSOLUTE_Y_STATE_0,
ORA_ABSOLUTE_Y_STATE_1,
ORA_ABSOLUTE_Y_STATE_2,
ORA_ABSOLUTE_Y_STATE_3,
ORA_ABSOLUTE_Y_STATE_4,
ORA_ABSOLUTE_Y_STATE_5,
ORA_ABSOLUTE_Y_STATE_6,
ORA_ABSOLUTE_Y_STATE_7,
ORA_ABSOLUTE_Y_STATE_8,
ORA_ABSOLUTE_Y_STATE_9,


ORA_IMMEDIATE_STATE_0,
ORA_IMMEDIATE_STATE_1,
ORA_IMMEDIATE_STATE_2,
ORA_IMMEDIATE_STATE_3,
ORA_IMMEDIATE_STATE_4,
ORA_IMMEDIATE_STATE_5,
ORA_IMMEDIATE_STATE_6,
ORA_IMMEDIATE_STATE_7,
ORA_IMMEDIATE_STATE_8,
ORA_IMMEDIATE_STATE_9,


ORA_INDIRECT_X_STATE_0,
ORA_INDIRECT_X_STATE_1,
ORA_INDIRECT_X_STATE_2,
ORA_INDIRECT_X_STATE_3,
ORA_INDIRECT_X_STATE_4,
ORA_INDIRECT_X_STATE_5,
ORA_INDIRECT_X_STATE_6,
ORA_INDIRECT_X_STATE_7,
ORA_INDIRECT_X_STATE_8,
ORA_INDIRECT_X_STATE_9,


ORA_INDIRECT_Y_STATE_0,
ORA_INDIRECT_Y_STATE_1,
ORA_INDIRECT_Y_STATE_2,
ORA_INDIRECT_Y_STATE_3,
ORA_INDIRECT_Y_STATE_4,
ORA_INDIRECT_Y_STATE_5,
ORA_INDIRECT_Y_STATE_6,
ORA_INDIRECT_Y_STATE_7,
ORA_INDIRECT_Y_STATE_8,
ORA_INDIRECT_Y_STATE_9,


ORA_ZERO_PAGE_STATE_0,
ORA_ZERO_PAGE_STATE_1,
ORA_ZERO_PAGE_STATE_2,
ORA_ZERO_PAGE_STATE_3,
ORA_ZERO_PAGE_STATE_4,
ORA_ZERO_PAGE_STATE_5,
ORA_ZERO_PAGE_STATE_6,
ORA_ZERO_PAGE_STATE_7,
ORA_ZERO_PAGE_STATE_8,
ORA_ZERO_PAGE_STATE_9,


ORA_ZERO_PAGE_X_STATE_0,
ORA_ZERO_PAGE_X_STATE_1,
ORA_ZERO_PAGE_X_STATE_2,
ORA_ZERO_PAGE_X_STATE_3,
ORA_ZERO_PAGE_X_STATE_4,
ORA_ZERO_PAGE_X_STATE_5,
ORA_ZERO_PAGE_X_STATE_6,
ORA_ZERO_PAGE_X_STATE_7,
ORA_ZERO_PAGE_X_STATE_8,
ORA_ZERO_PAGE_X_STATE_9,


PHA_IMPLIED_STATE_0,
PHA_IMPLIED_STATE_1,
PHA_IMPLIED_STATE_2,
PHA_IMPLIED_STATE_3,
PHA_IMPLIED_STATE_4,
PHA_IMPLIED_STATE_5,
PHA_IMPLIED_STATE_6,
PHA_IMPLIED_STATE_7,
PHA_IMPLIED_STATE_8,
PHA_IMPLIED_STATE_9,


PHP_IMPLIED_STATE_0,
PHP_IMPLIED_STATE_1,
PHP_IMPLIED_STATE_2,
PHP_IMPLIED_STATE_3,
PHP_IMPLIED_STATE_4,
PHP_IMPLIED_STATE_5,
PHP_IMPLIED_STATE_6,
PHP_IMPLIED_STATE_7,
PHP_IMPLIED_STATE_8,
PHP_IMPLIED_STATE_9,


PLA_IMPLIED_STATE_0,
PLA_IMPLIED_STATE_1,
PLA_IMPLIED_STATE_2,
PLA_IMPLIED_STATE_3,
PLA_IMPLIED_STATE_4,
PLA_IMPLIED_STATE_5,
PLA_IMPLIED_STATE_6,
PLA_IMPLIED_STATE_7,
PLA_IMPLIED_STATE_8,
PLA_IMPLIED_STATE_9,


PLP_IMPLIED_STATE_0,
PLP_IMPLIED_STATE_1,
PLP_IMPLIED_STATE_2,
PLP_IMPLIED_STATE_3,
PLP_IMPLIED_STATE_4,
PLP_IMPLIED_STATE_5,
PLP_IMPLIED_STATE_6,
PLP_IMPLIED_STATE_7,
PLP_IMPLIED_STATE_8,
PLP_IMPLIED_STATE_9,


RESET_INTERNAL_STATE_0,
RESET_INTERNAL_STATE_1,
RESET_INTERNAL_STATE_2,
RESET_INTERNAL_STATE_3,
RESET_INTERNAL_STATE_4,
RESET_INTERNAL_STATE_5,
RESET_INTERNAL_STATE_6,
RESET_INTERNAL_STATE_7,
RESET_INTERNAL_STATE_8,
RESET_INTERNAL_STATE_9,


ROL_ABSOLUTE_STATE_0,
ROL_ABSOLUTE_STATE_1,
ROL_ABSOLUTE_STATE_2,
ROL_ABSOLUTE_STATE_3,
ROL_ABSOLUTE_STATE_4,
ROL_ABSOLUTE_STATE_5,
ROL_ABSOLUTE_STATE_6,
ROL_ABSOLUTE_STATE_7,
ROL_ABSOLUTE_STATE_8,
ROL_ABSOLUTE_STATE_9,


ROL_ABSOLUTE_X_STATE_0,
ROL_ABSOLUTE_X_STATE_1,
ROL_ABSOLUTE_X_STATE_2,
ROL_ABSOLUTE_X_STATE_3,
ROL_ABSOLUTE_X_STATE_4,
ROL_ABSOLUTE_X_STATE_5,
ROL_ABSOLUTE_X_STATE_6,
ROL_ABSOLUTE_X_STATE_7,
ROL_ABSOLUTE_X_STATE_8,
ROL_ABSOLUTE_X_STATE_9,


ROL_ACCUMULATOR_STATE_0,
ROL_ACCUMULATOR_STATE_1,
ROL_ACCUMULATOR_STATE_2,
ROL_ACCUMULATOR_STATE_3,
ROL_ACCUMULATOR_STATE_4,
ROL_ACCUMULATOR_STATE_5,
ROL_ACCUMULATOR_STATE_6,
ROL_ACCUMULATOR_STATE_7,
ROL_ACCUMULATOR_STATE_8,
ROL_ACCUMULATOR_STATE_9,


ROL_ZERO_PAGE_STATE_0,
ROL_ZERO_PAGE_STATE_1,
ROL_ZERO_PAGE_STATE_2,
ROL_ZERO_PAGE_STATE_3,
ROL_ZERO_PAGE_STATE_4,
ROL_ZERO_PAGE_STATE_5,
ROL_ZERO_PAGE_STATE_6,
ROL_ZERO_PAGE_STATE_7,
ROL_ZERO_PAGE_STATE_8,
ROL_ZERO_PAGE_STATE_9,


ROL_ZERO_PAGE_X_STATE_0,
ROL_ZERO_PAGE_X_STATE_1,
ROL_ZERO_PAGE_X_STATE_2,
ROL_ZERO_PAGE_X_STATE_3,
ROL_ZERO_PAGE_X_STATE_4,
ROL_ZERO_PAGE_X_STATE_5,
ROL_ZERO_PAGE_X_STATE_6,
ROL_ZERO_PAGE_X_STATE_7,
ROL_ZERO_PAGE_X_STATE_8,
ROL_ZERO_PAGE_X_STATE_9,


ROR_ABSOLUTE_STATE_0,
ROR_ABSOLUTE_STATE_1,
ROR_ABSOLUTE_STATE_2,
ROR_ABSOLUTE_STATE_3,
ROR_ABSOLUTE_STATE_4,
ROR_ABSOLUTE_STATE_5,
ROR_ABSOLUTE_STATE_6,
ROR_ABSOLUTE_STATE_7,
ROR_ABSOLUTE_STATE_8,
ROR_ABSOLUTE_STATE_9,


ROR_ABSOLUTE_X_STATE_0,
ROR_ABSOLUTE_X_STATE_1,
ROR_ABSOLUTE_X_STATE_2,
ROR_ABSOLUTE_X_STATE_3,
ROR_ABSOLUTE_X_STATE_4,
ROR_ABSOLUTE_X_STATE_5,
ROR_ABSOLUTE_X_STATE_6,
ROR_ABSOLUTE_X_STATE_7,
ROR_ABSOLUTE_X_STATE_8,
ROR_ABSOLUTE_X_STATE_9,


ROR_ACCUMULATOR_STATE_0,
ROR_ACCUMULATOR_STATE_1,
ROR_ACCUMULATOR_STATE_2,
ROR_ACCUMULATOR_STATE_3,
ROR_ACCUMULATOR_STATE_4,
ROR_ACCUMULATOR_STATE_5,
ROR_ACCUMULATOR_STATE_6,
ROR_ACCUMULATOR_STATE_7,
ROR_ACCUMULATOR_STATE_8,
ROR_ACCUMULATOR_STATE_9,


ROR_ZERO_PAGE_STATE_0,
ROR_ZERO_PAGE_STATE_1,
ROR_ZERO_PAGE_STATE_2,
ROR_ZERO_PAGE_STATE_3,
ROR_ZERO_PAGE_STATE_4,
ROR_ZERO_PAGE_STATE_5,
ROR_ZERO_PAGE_STATE_6,
ROR_ZERO_PAGE_STATE_7,
ROR_ZERO_PAGE_STATE_8,
ROR_ZERO_PAGE_STATE_9,


ROR_ZERO_PAGE_X_STATE_0,
ROR_ZERO_PAGE_X_STATE_1,
ROR_ZERO_PAGE_X_STATE_2,
ROR_ZERO_PAGE_X_STATE_3,
ROR_ZERO_PAGE_X_STATE_4,
ROR_ZERO_PAGE_X_STATE_5,
ROR_ZERO_PAGE_X_STATE_6,
ROR_ZERO_PAGE_X_STATE_7,
ROR_ZERO_PAGE_X_STATE_8,
ROR_ZERO_PAGE_X_STATE_9,


RTI_IMPLIED_STATE_0,
RTI_IMPLIED_STATE_1,
RTI_IMPLIED_STATE_2,
RTI_IMPLIED_STATE_3,
RTI_IMPLIED_STATE_4,
RTI_IMPLIED_STATE_5,
RTI_IMPLIED_STATE_6,
RTI_IMPLIED_STATE_7,
RTI_IMPLIED_STATE_8,
RTI_IMPLIED_STATE_9,


RTS_IMPLIED_STATE_0,
RTS_IMPLIED_STATE_1,
RTS_IMPLIED_STATE_2,
RTS_IMPLIED_STATE_3,
RTS_IMPLIED_STATE_4,
RTS_IMPLIED_STATE_5,
RTS_IMPLIED_STATE_6,
RTS_IMPLIED_STATE_7,
RTS_IMPLIED_STATE_8,
RTS_IMPLIED_STATE_9,


SBC_ABSOLUTE_STATE_0,
SBC_ABSOLUTE_STATE_1,
SBC_ABSOLUTE_STATE_2,
SBC_ABSOLUTE_STATE_3,
SBC_ABSOLUTE_STATE_4,
SBC_ABSOLUTE_STATE_5,
SBC_ABSOLUTE_STATE_6,
SBC_ABSOLUTE_STATE_7,
SBC_ABSOLUTE_STATE_8,
SBC_ABSOLUTE_STATE_9,


SBC_ABSOLUTE_X_STATE_0,
SBC_ABSOLUTE_X_STATE_1,
SBC_ABSOLUTE_X_STATE_2,
SBC_ABSOLUTE_X_STATE_3,
SBC_ABSOLUTE_X_STATE_4,
SBC_ABSOLUTE_X_STATE_5,
SBC_ABSOLUTE_X_STATE_6,
SBC_ABSOLUTE_X_STATE_7,
SBC_ABSOLUTE_X_STATE_8,
SBC_ABSOLUTE_X_STATE_9,


SBC_ABSOLUTE_Y_STATE_0,
SBC_ABSOLUTE_Y_STATE_1,
SBC_ABSOLUTE_Y_STATE_2,
SBC_ABSOLUTE_Y_STATE_3,
SBC_ABSOLUTE_Y_STATE_4,
SBC_ABSOLUTE_Y_STATE_5,
SBC_ABSOLUTE_Y_STATE_6,
SBC_ABSOLUTE_Y_STATE_7,
SBC_ABSOLUTE_Y_STATE_8,
SBC_ABSOLUTE_Y_STATE_9,


SBC_IMMEDIATE_STATE_0,
SBC_IMMEDIATE_STATE_1,
SBC_IMMEDIATE_STATE_2,
SBC_IMMEDIATE_STATE_3,
SBC_IMMEDIATE_STATE_4,
SBC_IMMEDIATE_STATE_5,
SBC_IMMEDIATE_STATE_6,
SBC_IMMEDIATE_STATE_7,
SBC_IMMEDIATE_STATE_8,
SBC_IMMEDIATE_STATE_9,


SBC_INDIRECT_X_STATE_0,
SBC_INDIRECT_X_STATE_1,
SBC_INDIRECT_X_STATE_2,
SBC_INDIRECT_X_STATE_3,
SBC_INDIRECT_X_STATE_4,
SBC_INDIRECT_X_STATE_5,
SBC_INDIRECT_X_STATE_6,
SBC_INDIRECT_X_STATE_7,
SBC_INDIRECT_X_STATE_8,
SBC_INDIRECT_X_STATE_9,


SBC_INDIRECT_Y_STATE_0,
SBC_INDIRECT_Y_STATE_1,
SBC_INDIRECT_Y_STATE_2,
SBC_INDIRECT_Y_STATE_3,
SBC_INDIRECT_Y_STATE_4,
SBC_INDIRECT_Y_STATE_5,
SBC_INDIRECT_Y_STATE_6,
SBC_INDIRECT_Y_STATE_7,
SBC_INDIRECT_Y_STATE_8,
SBC_INDIRECT_Y_STATE_9,


SBC_ZERO_PAGE_STATE_0,
SBC_ZERO_PAGE_STATE_1,
SBC_ZERO_PAGE_STATE_2,
SBC_ZERO_PAGE_STATE_3,
SBC_ZERO_PAGE_STATE_4,
SBC_ZERO_PAGE_STATE_5,
SBC_ZERO_PAGE_STATE_6,
SBC_ZERO_PAGE_STATE_7,
SBC_ZERO_PAGE_STATE_8,
SBC_ZERO_PAGE_STATE_9,


SBC_ZERO_PAGE_X_STATE_0,
SBC_ZERO_PAGE_X_STATE_1,
SBC_ZERO_PAGE_X_STATE_2,
SBC_ZERO_PAGE_X_STATE_3,
SBC_ZERO_PAGE_X_STATE_4,
SBC_ZERO_PAGE_X_STATE_5,
SBC_ZERO_PAGE_X_STATE_6,
SBC_ZERO_PAGE_X_STATE_7,
SBC_ZERO_PAGE_X_STATE_8,
SBC_ZERO_PAGE_X_STATE_9,


SEC_IMPLIED_STATE_0,
SEC_IMPLIED_STATE_1,
SEC_IMPLIED_STATE_2,
SEC_IMPLIED_STATE_3,
SEC_IMPLIED_STATE_4,
SEC_IMPLIED_STATE_5,
SEC_IMPLIED_STATE_6,
SEC_IMPLIED_STATE_7,
SEC_IMPLIED_STATE_8,
SEC_IMPLIED_STATE_9,


SED_IMPLIED_STATE_0,
SED_IMPLIED_STATE_1,
SED_IMPLIED_STATE_2,
SED_IMPLIED_STATE_3,
SED_IMPLIED_STATE_4,
SED_IMPLIED_STATE_5,
SED_IMPLIED_STATE_6,
SED_IMPLIED_STATE_7,
SED_IMPLIED_STATE_8,
SED_IMPLIED_STATE_9,


SEI_IMPLIED_STATE_0,
SEI_IMPLIED_STATE_1,
SEI_IMPLIED_STATE_2,
SEI_IMPLIED_STATE_3,
SEI_IMPLIED_STATE_4,
SEI_IMPLIED_STATE_5,
SEI_IMPLIED_STATE_6,
SEI_IMPLIED_STATE_7,
SEI_IMPLIED_STATE_8,
SEI_IMPLIED_STATE_9,


STA_ABSOLUTE_STATE_0,
STA_ABSOLUTE_STATE_1,
STA_ABSOLUTE_STATE_2,
STA_ABSOLUTE_STATE_3,
STA_ABSOLUTE_STATE_4,
STA_ABSOLUTE_STATE_5,
STA_ABSOLUTE_STATE_6,
STA_ABSOLUTE_STATE_7,
STA_ABSOLUTE_STATE_8,
STA_ABSOLUTE_STATE_9,


STA_ABSOLUTE_Y_STATE_0,
STA_ABSOLUTE_Y_STATE_1,
STA_ABSOLUTE_Y_STATE_2,
STA_ABSOLUTE_Y_STATE_3,
STA_ABSOLUTE_Y_STATE_4,
STA_ABSOLUTE_Y_STATE_5,
STA_ABSOLUTE_Y_STATE_6,
STA_ABSOLUTE_Y_STATE_7,
STA_ABSOLUTE_Y_STATE_8,
STA_ABSOLUTE_Y_STATE_9,


STA_INDIRECT_X_STATE_0,
STA_INDIRECT_X_STATE_1,
STA_INDIRECT_X_STATE_2,
STA_INDIRECT_X_STATE_3,
STA_INDIRECT_X_STATE_4,
STA_INDIRECT_X_STATE_5,
STA_INDIRECT_X_STATE_6,
STA_INDIRECT_X_STATE_7,
STA_INDIRECT_X_STATE_8,
STA_INDIRECT_X_STATE_9,


STA_INDIRECT_Y_STATE_0,
STA_INDIRECT_Y_STATE_1,
STA_INDIRECT_Y_STATE_2,
STA_INDIRECT_Y_STATE_3,
STA_INDIRECT_Y_STATE_4,
STA_INDIRECT_Y_STATE_5,
STA_INDIRECT_Y_STATE_6,
STA_INDIRECT_Y_STATE_7,
STA_INDIRECT_Y_STATE_8,
STA_INDIRECT_Y_STATE_9,


STA_ZERO_PAGE_STATE_0,
STA_ZERO_PAGE_STATE_1,
STA_ZERO_PAGE_STATE_2,
STA_ZERO_PAGE_STATE_3,
STA_ZERO_PAGE_STATE_4,
STA_ZERO_PAGE_STATE_5,
STA_ZERO_PAGE_STATE_6,
STA_ZERO_PAGE_STATE_7,
STA_ZERO_PAGE_STATE_8,
STA_ZERO_PAGE_STATE_9,


STA_ZERO_PAGE_X_STATE_0,
STA_ZERO_PAGE_X_STATE_1,
STA_ZERO_PAGE_X_STATE_2,
STA_ZERO_PAGE_X_STATE_3,
STA_ZERO_PAGE_X_STATE_4,
STA_ZERO_PAGE_X_STATE_5,
STA_ZERO_PAGE_X_STATE_6,
STA_ZERO_PAGE_X_STATE_7,
STA_ZERO_PAGE_X_STATE_8,
STA_ZERO_PAGE_X_STATE_9,


STA_ABSOLUTE_X_STATE_0,
STA_ABSOLUTE_X_STATE_1,
STA_ABSOLUTE_X_STATE_2,
STA_ABSOLUTE_X_STATE_3,
STA_ABSOLUTE_X_STATE_4,
STA_ABSOLUTE_X_STATE_5,
STA_ABSOLUTE_X_STATE_6,
STA_ABSOLUTE_X_STATE_7,
STA_ABSOLUTE_X_STATE_8,
STA_ABSOLUTE_X_STATE_9,


S_IRQ_INTERNAL_STATE_0,
S_IRQ_INTERNAL_STATE_1,
S_IRQ_INTERNAL_STATE_2,
S_IRQ_INTERNAL_STATE_3,
S_IRQ_INTERNAL_STATE_4,
S_IRQ_INTERNAL_STATE_5,
S_IRQ_INTERNAL_STATE_6,
S_IRQ_INTERNAL_STATE_7,
S_IRQ_INTERNAL_STATE_8,
S_IRQ_INTERNAL_STATE_9,


S_NMI_INTERNAL_STATE_0,
S_NMI_INTERNAL_STATE_1,
S_NMI_INTERNAL_STATE_2,
S_NMI_INTERNAL_STATE_3,
S_NMI_INTERNAL_STATE_4,
S_NMI_INTERNAL_STATE_5,
S_NMI_INTERNAL_STATE_6,
S_NMI_INTERNAL_STATE_7,
S_NMI_INTERNAL_STATE_8,
S_NMI_INTERNAL_STATE_9,


STX_ABSOLUTE_STATE_0,
STX_ABSOLUTE_STATE_1,
STX_ABSOLUTE_STATE_2,
STX_ABSOLUTE_STATE_3,
STX_ABSOLUTE_STATE_4,
STX_ABSOLUTE_STATE_5,
STX_ABSOLUTE_STATE_6,
STX_ABSOLUTE_STATE_7,
STX_ABSOLUTE_STATE_8,
STX_ABSOLUTE_STATE_9,


STX_ZERO_PAGE_STATE_0,
STX_ZERO_PAGE_STATE_1,
STX_ZERO_PAGE_STATE_2,
STX_ZERO_PAGE_STATE_3,
STX_ZERO_PAGE_STATE_4,
STX_ZERO_PAGE_STATE_5,
STX_ZERO_PAGE_STATE_6,
STX_ZERO_PAGE_STATE_7,
STX_ZERO_PAGE_STATE_8,
STX_ZERO_PAGE_STATE_9,


STX_ZERO_PAGE_Y_STATE_0,
STX_ZERO_PAGE_Y_STATE_1,
STX_ZERO_PAGE_Y_STATE_2,
STX_ZERO_PAGE_Y_STATE_3,
STX_ZERO_PAGE_Y_STATE_4,
STX_ZERO_PAGE_Y_STATE_5,
STX_ZERO_PAGE_Y_STATE_6,
STX_ZERO_PAGE_Y_STATE_7,
STX_ZERO_PAGE_Y_STATE_8,
STX_ZERO_PAGE_Y_STATE_9,


STY_ABSOLUTE_STATE_0,
STY_ABSOLUTE_STATE_1,
STY_ABSOLUTE_STATE_2,
STY_ABSOLUTE_STATE_3,
STY_ABSOLUTE_STATE_4,
STY_ABSOLUTE_STATE_5,
STY_ABSOLUTE_STATE_6,
STY_ABSOLUTE_STATE_7,
STY_ABSOLUTE_STATE_8,
STY_ABSOLUTE_STATE_9,


STY_ZERO_PAGE_STATE_0,
STY_ZERO_PAGE_STATE_1,
STY_ZERO_PAGE_STATE_2,
STY_ZERO_PAGE_STATE_3,
STY_ZERO_PAGE_STATE_4,
STY_ZERO_PAGE_STATE_5,
STY_ZERO_PAGE_STATE_6,
STY_ZERO_PAGE_STATE_7,
STY_ZERO_PAGE_STATE_8,
STY_ZERO_PAGE_STATE_9,


STY_ZERO_PAGE_X_STATE_0,
STY_ZERO_PAGE_X_STATE_1,
STY_ZERO_PAGE_X_STATE_2,
STY_ZERO_PAGE_X_STATE_3,
STY_ZERO_PAGE_X_STATE_4,
STY_ZERO_PAGE_X_STATE_5,
STY_ZERO_PAGE_X_STATE_6,
STY_ZERO_PAGE_X_STATE_7,
STY_ZERO_PAGE_X_STATE_8,
STY_ZERO_PAGE_X_STATE_9,


TAX_IMPLIED_STATE_0,
TAX_IMPLIED_STATE_1,
TAX_IMPLIED_STATE_2,
TAX_IMPLIED_STATE_3,
TAX_IMPLIED_STATE_4,
TAX_IMPLIED_STATE_5,
TAX_IMPLIED_STATE_6,
TAX_IMPLIED_STATE_7,
TAX_IMPLIED_STATE_8,
TAX_IMPLIED_STATE_9,


TAY_IMPLIED_STATE_0,
TAY_IMPLIED_STATE_1,
TAY_IMPLIED_STATE_2,
TAY_IMPLIED_STATE_3,
TAY_IMPLIED_STATE_4,
TAY_IMPLIED_STATE_5,
TAY_IMPLIED_STATE_6,
TAY_IMPLIED_STATE_7,
TAY_IMPLIED_STATE_8,
TAY_IMPLIED_STATE_9,


TSX_IMPLIED_STATE_0,
TSX_IMPLIED_STATE_1,
TSX_IMPLIED_STATE_2,
TSX_IMPLIED_STATE_3,
TSX_IMPLIED_STATE_4,
TSX_IMPLIED_STATE_5,
TSX_IMPLIED_STATE_6,
TSX_IMPLIED_STATE_7,
TSX_IMPLIED_STATE_8,
TSX_IMPLIED_STATE_9,


TXA_IMPLIED_STATE_0,
TXA_IMPLIED_STATE_1,
TXA_IMPLIED_STATE_2,
TXA_IMPLIED_STATE_3,
TXA_IMPLIED_STATE_4,
TXA_IMPLIED_STATE_5,
TXA_IMPLIED_STATE_6,
TXA_IMPLIED_STATE_7,
TXA_IMPLIED_STATE_8,
TXA_IMPLIED_STATE_9,


TXS_IMPLIED_STATE_0,
TXS_IMPLIED_STATE_1,
TXS_IMPLIED_STATE_2,
TXS_IMPLIED_STATE_3,
TXS_IMPLIED_STATE_4,
TXS_IMPLIED_STATE_5,
TXS_IMPLIED_STATE_6,
TXS_IMPLIED_STATE_7,
TXS_IMPLIED_STATE_8,
TXS_IMPLIED_STATE_9,


--- end generated code




	HOSED,
NEW_INSTRUCTION,
FETCH_0,
FETCH_INSTRUCTION,

ABSOLUTE_0,
ABSOLUTE_1,
ABSOLUTE_2,
ABSOLUTE_3,
ABSOLUTE_4,
ABSOLUTE_5,


ABSOLUTE_X_0,


ABSOLUTE_Y_0,



IMMEDIATE_0,
IMMEDIATE_1,
IMMEDIATE_2,



INDIRECT_X_0,



INDIRECT_Y_0,



ZERO_PAGE_0,



ZERO_PAGE_X_0,


ZERO_PAGE_Y_0,


RELATIVE_0,


IMPLIED_0,


ACCUMULATOR_0,


INDIRECT_0,


INTERNAL_0,

LDX_IMMEDIATE_0,
LDY_IMMEDIATE_0,
LDA_IMMEDIATE_0


);



constant LO:     std_logic:='0';
constant HI:     std_logic:='1';
constant ADC_ABSOLUTE     : std_logic_vector (7 downto 0):=  "01101101";
constant ADC_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "01111101";
constant ADC_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "01111001";
constant ADC_IMMEDIATE    : std_logic_vector (7 downto 0):=  "01101001";
constant ADC_INDIRECT_X   : std_logic_vector (7 downto 0):=  "01100001";
constant ADC_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "01110001";
constant ADC_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "01100101";
constant ADC_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "01110101";
constant AND_ABSOLUTE     : std_logic_vector (7 downto 0):=  "00101101";
constant AND_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "00111101";
constant AND_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "00111001";
constant AND_IMMEDIATE    : std_logic_vector (7 downto 0):=  "00101001";
constant AND_INDIRECT_X   : std_logic_vector (7 downto 0):=  "00100001";
constant AND_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "00110001";
constant AND_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "00100101";
constant AND_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "00110101";
constant ASL_ABSOLUTE     : std_logic_vector (7 downto 0):=  "00001110";
constant ASL_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "00011110";
constant ASL_ACCUMULATOR  : std_logic_vector (7 downto 0):=  "00001010";
constant ASL_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "00000110";
constant ASL_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "00010110";
constant BCC_RELATIVE     : std_logic_vector (7 downto 0):=  "10010000";
constant BCS_RELATIVE     : std_logic_vector (7 downto 0):=  "10110000";
constant BEQ_RELATIVE     : std_logic_vector (7 downto 0):=  "11110000";
constant BIT_ABSOLUTE     : std_logic_vector (7 downto 0):=  "00101100";
constant BIT_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "00100100";
constant BMI_RELATIVE     : std_logic_vector (7 downto 0):=  "00110000";
constant BNE_RELATIVE     : std_logic_vector (7 downto 0):=  "11010000";
constant BPL_RELATIVE     : std_logic_vector (7 downto 0):=  "00010000";
constant BRK_IMPLIED      : std_logic_vector (7 downto 0):=  "00000000";
constant BVC_RELATIVE     : std_logic_vector (7 downto 0):=  "01010000";
constant BVS_RELATIVE     : std_logic_vector (7 downto 0):=  "01110000";
constant CLC_IMPLIED      : std_logic_vector (7 downto 0):=  "00011000";
constant CLD_IMPLIED      : std_logic_vector (7 downto 0):=  "11011000";
constant CLI_IMPLIED      : std_logic_vector (7 downto 0):=  "01011000";
constant CLV_IMPLIED      : std_logic_vector (7 downto 0):=  "10111000";
constant CMP_ABSOLUTE     : std_logic_vector (7 downto 0):=  "11001101";
constant CMP_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "11011101";
constant CMP_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "11011001";
constant CMP_IMMEDIATE    : std_logic_vector (7 downto 0):=  "11001001";
constant CMP_INDIRECT_X   : std_logic_vector (7 downto 0):=  "11000001";
constant CMP_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "11010001";
constant CMP_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "11000101";
constant CMP_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "11010101";
constant CPX_ABSOLUTE     : std_logic_vector (7 downto 0):=  "11101100";
constant CPX_IMMEDIATE    : std_logic_vector (7 downto 0):=  "11100000";
constant CPX_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "11100100";
constant CPY_ABSOLUTE     : std_logic_vector (7 downto 0):=  "11001100";
constant CPY_IMMEDIATE    : std_logic_vector (7 downto 0):=  "11000000";
constant CPY_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "11000100";
constant DEC_ABSOLUTE     : std_logic_vector (7 downto 0):=  "11001110";
constant DEC_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "11011110";
constant DEC_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "11000110";
constant DEC_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "11010110";
constant DEX_IMPLIED      : std_logic_vector (7 downto 0):=  "11001010";
constant DEY_IMPLIED      : std_logic_vector (7 downto 0):=  "10001000";
constant EOR_ABSOLUTE     : std_logic_vector (7 downto 0):=  "01001101";
constant EOR_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "01011101";
constant EOR_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "01011001";
constant EOR_IMMEDIATE    : std_logic_vector (7 downto 0):=  "01001001";
constant EOR_INDIRECT_X   : std_logic_vector (7 downto 0):=  "01000001";
constant EOR_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "01010001";
constant EOR_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "01000101";
constant EOR_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "01010101";
constant INC_ABSOLUTE     : std_logic_vector (7 downto 0):=  "11101110";
constant INC_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "11111110";
constant INC_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "11100110";
constant INC_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "11110110";
constant INX_IMPLIED      : std_logic_vector (7 downto 0):=  "11101000";
constant INY_IMPLIED      : std_logic_vector (7 downto 0):=  "11001000";
constant JMP_ABSOLUTE     : std_logic_vector (7 downto 0):=  "01001100";
constant JMP_INDIRECT     : std_logic_vector (7 downto 0):=  "01101100";
constant JSR_ABSOLUTE     : std_logic_vector (7 downto 0):=  "00100000";
constant LDA_ABSOLUTE     : std_logic_vector (7 downto 0):=  "10101101";
constant LDA_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "10111101";
constant LDA_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "10111001";
constant LDA_IMMEDIATE    : std_logic_vector (7 downto 0):=  "10101001";
constant LDA_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "10100101";
constant LDA_INDIRECT_X   : std_logic_vector (7 downto 0):=  "10100001";
constant LDA_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "10110001";
constant LDA_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "10110101";
constant LDX_ABSOLUTE     : std_logic_vector (7 downto 0):=  "10101110";
constant LDX_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "10111110";
constant LDX_IMMEDIATE    : std_logic_vector (7 downto 0):=  "10100010";
constant LDX_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "10100110";
constant LDX_ZERO_PAGE_Y  : std_logic_vector (7 downto 0):=  "10110110";
constant LDY_ABSOLUTE     : std_logic_vector (7 downto 0):=  "10101100";
constant LDY_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "10111100";
constant LDY_IMMEDIATE    : std_logic_vector (7 downto 0):=  "10100000";
constant LDY_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "10100100";
constant LDY_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "10110100";
constant LSR_ABSOLUTE     : std_logic_vector (7 downto 0):=  "01001110";
constant LSR_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "01011110";
constant LSR_ACCUMULATOR  : std_logic_vector (7 downto 0):=  "01001010";
constant LSR_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "01000110";
constant LSR_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "01010110";
constant NOP_IMPLIED      : std_logic_vector (7 downto 0):=  "11101010";
constant ORA_ABSOLUTE     : std_logic_vector (7 downto 0):=  "00001101";
constant ORA_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "00011101";
constant ORA_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "00011001";
constant ORA_IMMEDIATE    : std_logic_vector (7 downto 0):=  "00001001";
constant ORA_INDIRECT_X   : std_logic_vector (7 downto 0):=  "00000001";
constant ORA_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "00010001";
constant ORA_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "00000101";
constant ORA_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "00010101";
constant PHA_IMPLIED      : std_logic_vector (7 downto 0):=  "01001000";
constant PHP_IMPLIED      : std_logic_vector (7 downto 0):=  "00001000";
constant PLA_IMPLIED      : std_logic_vector (7 downto 0):=  "01101000";
constant PLP_IMPLIED      : std_logic_vector (7 downto 0):=  "00101000";
constant RESET_INTERNAL   : std_logic_vector (7 downto 0):=  "00000011";
constant ROL_ABSOLUTE     : std_logic_vector (7 downto 0):=  "00101110";
constant ROL_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "00111110";
constant ROL_ACCUMULATOR  : std_logic_vector (7 downto 0):=  "00101010";
constant ROL_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "00100110";
constant ROL_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "00110110";
constant ROR_ABSOLUTE     : std_logic_vector (7 downto 0):=  "01101110";
constant ROR_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "01111110";
constant ROR_ACCUMULATOR  : std_logic_vector (7 downto 0):=  "01101010";
constant ROR_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "01100110";
constant ROR_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "01110110";
constant RTI_IMPLIED      : std_logic_vector (7 downto 0):=  "01000000";
constant RTS_IMPLIED      : std_logic_vector (7 downto 0):=  "01100000";
constant SBC_ABSOLUTE     : std_logic_vector (7 downto 0):=  "11101101";
constant SBC_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "11111101";
constant SBC_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "11111001";
constant SBC_IMMEDIATE    : std_logic_vector (7 downto 0):=  "11101001";
constant SBC_INDIRECT_X   : std_logic_vector (7 downto 0):=  "11100001";
constant SBC_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "11110001";
constant SBC_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "11100101";
constant SBC_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "11110101";
constant SEC_IMPLIED      : std_logic_vector (7 downto 0):=  "00111000";
constant SED_IMPLIED      : std_logic_vector (7 downto 0):=  "11111000";
constant SEI_IMPLIED      : std_logic_vector (7 downto 0):=  "01111000";
constant STA_ABSOLUTE     : std_logic_vector (7 downto 0):=  "10001101";
constant STA_ABSOLUTE_Y   : std_logic_vector (7 downto 0):=  "10011001";
constant STA_INDIRECT_X   : std_logic_vector (7 downto 0):=  "10000001";
constant STA_INDIRECT_Y   : std_logic_vector (7 downto 0):=  "10010001";
constant STA_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "10000101";
constant STA_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "10010101";
constant STA_ABSOLUTE_X   : std_logic_vector (7 downto 0):=  "10011101";
constant S_IRQ_INTERNAL   : std_logic_vector (7 downto 0):=  "01000011";
constant S_NMI_INTERNAL   : std_logic_vector (7 downto 0):=  "00110011";
constant STX_ABSOLUTE     : std_logic_vector (7 downto 0):=  "10001110";
constant STX_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "10000110";
constant STX_ZERO_PAGE_Y  : std_logic_vector (7 downto 0):=  "10010110";
constant STY_ABSOLUTE     : std_logic_vector (7 downto 0):=  "10001100";
constant STY_ZERO_PAGE    : std_logic_vector (7 downto 0):=  "10000100";
constant STY_ZERO_PAGE_X  : std_logic_vector (7 downto 0):=  "10010100";
constant TAX_IMPLIED      : std_logic_vector (7 downto 0):=  "10101010";
constant TAY_IMPLIED      : std_logic_vector (7 downto 0):=  "10101000";
constant TSX_IMPLIED      : std_logic_vector (7 downto 0):=  "10111010";
constant TXA_IMPLIED      : std_logic_vector (7 downto 0):=  "10001010";
constant TXS_IMPLIED      : std_logic_vector (7 downto 0):=  "10011010";
constant TYA_IMPLIED      : std_logic_vector (7 downto 0):=  "10011000";

constant NO_WRITE_TO_MEM: std_logic:='1';
constant NO_READ_FROM_MEM: std_logic:='1';

signal mem_addr:  std_logic_vector(15 downto 0);
signal offset: std_logic_vector(7 downto 0);


signal mem_addr_r:  std_logic_vector(15 downto 0);
signal offset_r: std_logic_vector(7 downto 0);




signal current_state, next_state: machine_state;
signal byte_read: std_logic_vector(7 downto 0);

--- addressing modes
	--- case ABSOLUTE   -----
	--- case ABSOLUTE_X -----
	--- case ABSOLUTE_Y -----
	--- case IMMEDIATE  -----
	--- case INDIRECT_X -----
	--- case INDIRECT_Y -----
	--- case ZERO_PAGE  -----
	--- case ZERO_PAGE_X-----
	--- case ZERO_PAGE_Y-----
	--- case RELATIVE ---
	--- case IMPLIED ---
	--- case ACCUMULATOR-----
	--- case INDIRECT ---
	--- case INTERNAL ---
--- end addressing modes


--signal  bnbuf:  std_logic;

signal dummy: std_logic;

--- misc. signals

signal tmp_data_r: std_logic_vector(7 downto 0);
signal  ar_r: std_logic_vector(15 downto 0);
signal ac_r, instruction_r: std_logic_vector(7 downto 0);
signal pc_r: std_logic_vector(15 downto 0);
signal x_r, y_r: std_logic_vector(7 downto 0);
signal addr_lo_r, addr_hi_r: std_logic_vector(7 downto 0);

signal tmp_data: std_logic_vector(7 downto 0);
signal instruction: std_logic_vector(7 downto 0);
signal ar: std_logic_vector(15 downto 0);
signal ac,x,y: std_logic_vector(7 downto 0);
signal pc: std_logic_vector(15 downto 0);
signal addr_lo, addr_hi: std_logic_vector(7 downto 0);


-- initial pc should really be in the FFXX range
constant  initial_pc : std_logic_vector(15 downto 0):="0000000000001000";
signal counter: std_logic_vector(3 downto 0);

------------------------------------------------------------------------
-- Module Implementation
------------------------------------------------------------------------

begin


----U1:	IBUFG port map (I => btn, O => bnbuf);
---  sequential

process(clock, reset)
begin
if (reset='0') then
	counter<="0000";
	pc_r<=initial_pc; 
	ac_r<=(others=>'0');
	x_r<=(others=>'0');
	y_r<=(others=>'0');
elsif (clock'event and clock='1') then
	counter<=counter+1;
	ar_r<=ar; 
	pc_r<=pc;
        addr_lo_r<= addr_lo;
        addr_hi_r<= addr_hi;
	x_r<=x;
	y_r<=y;
	ac_r<=ac;
	tmp_data_r<=tmp_data;
end if;
end process;

--- combinational


peep <= ac_r;
address<= ar_r;


process(clock, current_state)
begin
case current_state is



when ADC_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ADC_ABSOLUTE_STATE_1;

when ADC_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ADC_ABSOLUTE_STATE_2;

when ADC_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=ADC_ABSOLUTE_STATE_3;

when ADC_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=ADC_ABSOLUTE_STATE_4;

when ADC_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=ADC_ABSOLUTE_STATE_5;

when ADC_ABSOLUTE_STATE_5=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when ADC_ABSOLUTE_X_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when ADC_ABSOLUTE_Y_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ADC_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=ADC_IMMEDIATE_STATE_1;
when ADC_IMMEDIATE_STATE_1=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when ADC_INDIRECT_X_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when ADC_INDIRECT_Y_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ADC_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ADC_ZERO_PAGE_STATE_1;

when ADC_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ADC_ZERO_PAGE_STATE_2;

when ADC_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=ADC_ZERO_PAGE_STATE_3;

when ADC_ZERO_PAGE_STATE_3=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when ADC_ZERO_PAGE_X_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=ac_r+data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when AND_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=AND_ABSOLUTE_STATE_1;

when AND_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=AND_ABSOLUTE_STATE_2;

when AND_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=AND_ABSOLUTE_STATE_3;

when AND_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=AND_ABSOLUTE_STATE_4;

when AND_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=AND_ABSOLUTE_STATE_5;

when AND_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when AND_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when AND_ABSOLUTE_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when AND_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=AND_IMMEDIATE_STATE_1;
when AND_IMMEDIATE_STATE_1=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when AND_INDIRECT_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when AND_INDIRECT_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when AND_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=AND_ZERO_PAGE_STATE_1;

when AND_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=AND_ZERO_PAGE_STATE_2;

when AND_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=AND_ZERO_PAGE_STATE_3;

when AND_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when AND_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ASL_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ASL_ABSOLUTE_STATE_1;

when ASL_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ASL_ABSOLUTE_STATE_2;

when ASL_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=ASL_ABSOLUTE_STATE_3;

when ASL_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=ASL_ABSOLUTE_STATE_4;

when ASL_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=ASL_ABSOLUTE_STATE_5;

when ASL_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when ASL_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- accumulator NOT IMPLEMENTED ----
when ASL_ACCUMULATOR_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ASL_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ASL_ZERO_PAGE_STATE_1;

when ASL_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ASL_ZERO_PAGE_STATE_2;

when ASL_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=ASL_ZERO_PAGE_STATE_3;

when ASL_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when ASL_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BCC_RELATIVE_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BCS_RELATIVE_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BEQ_RELATIVE_STATE_0=> --- OPERATION

-- start from strings--
     if(offset_r>0) then 
     pc<=pc_r+offset_r; 
     else 
     pc<=pc_r-offset_r; 
     end if;

-- end  start from strings--
    next_state<=NEW_INSTRUCTION;



when BIT_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=BIT_ABSOLUTE_STATE_1;

when BIT_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=BIT_ABSOLUTE_STATE_2;

when BIT_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=BIT_ABSOLUTE_STATE_3;

when BIT_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=BIT_ABSOLUTE_STATE_4;

when BIT_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=BIT_ABSOLUTE_STATE_5;

when BIT_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when BIT_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=BIT_ZERO_PAGE_STATE_1;

when BIT_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=BIT_ZERO_PAGE_STATE_2;

when BIT_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=BIT_ZERO_PAGE_STATE_3;

when BIT_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BMI_RELATIVE_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BNE_RELATIVE_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BPL_RELATIVE_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when BRK_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BVC_RELATIVE_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  relative NOT IMPLEMENTED ----
when BVS_RELATIVE_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when CLC_IMPLIED_STATE_0=> --- OPERATION

-- start from strings--
--- DONE

-- end  start from strings--
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when CLD_IMPLIED_STATE_0=> --- OPERATION

-- start from strings--
--- DONE

-- end  start from strings--
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when CLI_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when CLV_IMPLIED_STATE_0=> --- OPERATION

-- start from strings--
--- DONE

-- end  start from strings--
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CMP_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=CMP_ABSOLUTE_STATE_1;

when CMP_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=CMP_ABSOLUTE_STATE_2;

when CMP_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=CMP_ABSOLUTE_STATE_3;

when CMP_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=CMP_ABSOLUTE_STATE_4;

when CMP_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=CMP_ABSOLUTE_STATE_5;

when CMP_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when CMP_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when CMP_ABSOLUTE_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CMP_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=CMP_IMMEDIATE_STATE_1;
when CMP_IMMEDIATE_STATE_1=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when CMP_INDIRECT_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when CMP_INDIRECT_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CMP_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=CMP_ZERO_PAGE_STATE_1;

when CMP_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=CMP_ZERO_PAGE_STATE_2;

when CMP_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=CMP_ZERO_PAGE_STATE_3;

when CMP_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when CMP_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CPX_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=CPX_ABSOLUTE_STATE_1;

when CPX_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=CPX_ABSOLUTE_STATE_2;

when CPX_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=CPX_ABSOLUTE_STATE_3;

when CPX_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=CPX_ABSOLUTE_STATE_4;

when CPX_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=CPX_ABSOLUTE_STATE_5;

when CPX_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CPX_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=CPX_IMMEDIATE_STATE_1;
when CPX_IMMEDIATE_STATE_1=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CPX_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=CPX_ZERO_PAGE_STATE_1;

when CPX_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=CPX_ZERO_PAGE_STATE_2;

when CPX_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=CPX_ZERO_PAGE_STATE_3;

when CPX_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CPY_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=CPY_ABSOLUTE_STATE_1;

when CPY_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=CPY_ABSOLUTE_STATE_2;

when CPY_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=CPY_ABSOLUTE_STATE_3;

when CPY_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=CPY_ABSOLUTE_STATE_4;

when CPY_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=CPY_ABSOLUTE_STATE_5;

when CPY_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CPY_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=CPY_IMMEDIATE_STATE_1;
when CPY_IMMEDIATE_STATE_1=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when CPY_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=CPY_ZERO_PAGE_STATE_1;

when CPY_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=CPY_ZERO_PAGE_STATE_2;

when CPY_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=CPY_ZERO_PAGE_STATE_3;

when CPY_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when DEC_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=DEC_ABSOLUTE_STATE_1;

when DEC_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=DEC_ABSOLUTE_STATE_2;

when DEC_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=DEC_ABSOLUTE_STATE_3;

when DEC_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=DEC_ABSOLUTE_STATE_4;

when DEC_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=DEC_ABSOLUTE_STATE_5;

when DEC_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when DEC_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when DEC_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=DEC_ZERO_PAGE_STATE_1;

when DEC_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=DEC_ZERO_PAGE_STATE_2;

when DEC_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=DEC_ZERO_PAGE_STATE_3;

when DEC_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when DEC_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when DEX_IMPLIED_STATE_0=> --- OPERATION

-- start from strings--
   x<=x_r-1;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when DEY_IMPLIED_STATE_0=> --- OPERATION

-- start from strings--
   y<=y_r-1;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when EOR_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=EOR_ABSOLUTE_STATE_1;

when EOR_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=EOR_ABSOLUTE_STATE_2;

when EOR_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=EOR_ABSOLUTE_STATE_3;

when EOR_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=EOR_ABSOLUTE_STATE_4;

when EOR_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=EOR_ABSOLUTE_STATE_5;

when EOR_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when EOR_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when EOR_ABSOLUTE_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when EOR_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=EOR_IMMEDIATE_STATE_1;
when EOR_IMMEDIATE_STATE_1=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when EOR_INDIRECT_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when EOR_INDIRECT_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when EOR_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=EOR_ZERO_PAGE_STATE_1;

when EOR_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=EOR_ZERO_PAGE_STATE_2;

when EOR_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=EOR_ZERO_PAGE_STATE_3;

when EOR_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when EOR_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when INC_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=INC_ABSOLUTE_STATE_1;

when INC_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=INC_ABSOLUTE_STATE_2;

when INC_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=INC_ABSOLUTE_STATE_3;

when INC_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=INC_ABSOLUTE_STATE_4;

when INC_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=INC_ABSOLUTE_STATE_5;

when INC_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when INC_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when INC_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=INC_ZERO_PAGE_STATE_1;

when INC_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=INC_ZERO_PAGE_STATE_2;

when INC_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=INC_ZERO_PAGE_STATE_3;

when INC_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when INC_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when INX_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when INY_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when JMP_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=JMP_ABSOLUTE_STATE_1;

when JMP_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=JMP_ABSOLUTE_STATE_2;

when JMP_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=JMP_ABSOLUTE_STATE_3;

when JMP_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=JMP_ABSOLUTE_STATE_4;

when JMP_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=JMP_ABSOLUTE_STATE_5;

when JMP_ABSOLUTE_STATE_5=> --- OPERATION

-- start from strings--
    pc<=addr_hi_r & addr_lo_r;

-- end  start from strings--
    next_state<=NEW_INSTRUCTION;


---indirect NOT IMPLEMENTED ----
when JMP_INDIRECT_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;



when JSR_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=JSR_ABSOLUTE_STATE_1;

when JSR_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=JSR_ABSOLUTE_STATE_2;

when JSR_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=JSR_ABSOLUTE_STATE_3;

when JSR_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=JSR_ABSOLUTE_STATE_4;

when JSR_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=JSR_ABSOLUTE_STATE_5;

when JSR_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;



when LDA_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LDA_ABSOLUTE_STATE_1;

when LDA_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LDA_ABSOLUTE_STATE_2;

when LDA_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=LDA_ABSOLUTE_STATE_3;

when LDA_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=LDA_ABSOLUTE_STATE_4;

when LDA_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=LDA_ABSOLUTE_STATE_5;

when LDA_ABSOLUTE_STATE_5=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when LDA_ABSOLUTE_X_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when LDA_ABSOLUTE_Y_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDA_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=LDA_IMMEDIATE_STATE_1;
when LDA_IMMEDIATE_STATE_1=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDA_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LDA_ZERO_PAGE_STATE_1;

when LDA_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LDA_ZERO_PAGE_STATE_2;

when LDA_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=LDA_ZERO_PAGE_STATE_3;

when LDA_ZERO_PAGE_STATE_3=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when LDA_INDIRECT_X_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when LDA_INDIRECT_Y_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when LDA_ZERO_PAGE_X_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   ac<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDX_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LDX_ABSOLUTE_STATE_1;

when LDX_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LDX_ABSOLUTE_STATE_2;

when LDX_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=LDX_ABSOLUTE_STATE_3;

when LDX_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=LDX_ABSOLUTE_STATE_4;

when LDX_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=LDX_ABSOLUTE_STATE_5;

when LDX_ABSOLUTE_STATE_5=> --- OPERATION

-- start from strings--
    rd<=LO;
   x<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when LDX_ABSOLUTE_Y_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   x<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDX_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=LDX_IMMEDIATE_STATE_1;
when LDX_IMMEDIATE_STATE_1=> --- OPERATION

-- start from strings--
    rd<=LO;
   x<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDX_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LDX_ZERO_PAGE_STATE_1;

when LDX_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LDX_ZERO_PAGE_STATE_2;

when LDX_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=LDX_ZERO_PAGE_STATE_3;

when LDX_ZERO_PAGE_STATE_3=> --- OPERATION

-- start from strings--
    rd<=LO;
   x<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- zeropage_y NOT IMPLEMENTED ----
when LDX_ZERO_PAGE_Y_STATE_0=> --- OPERATION

-- start from strings--
    rd<=LO;
   x<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDY_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LDY_ABSOLUTE_STATE_1;

when LDY_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LDY_ABSOLUTE_STATE_2;

when LDY_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=LDY_ABSOLUTE_STATE_3;

when LDY_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=LDY_ABSOLUTE_STATE_4;

when LDY_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=LDY_ABSOLUTE_STATE_5;

when LDY_ABSOLUTE_STATE_5=> --- OPERATION

-- start from strings--
  rd<=LO;
   y<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when LDY_ABSOLUTE_X_STATE_0=> --- OPERATION

-- start from strings--
  rd<=LO;
   y<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDY_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=LDY_IMMEDIATE_STATE_1;
when LDY_IMMEDIATE_STATE_1=> --- OPERATION

-- start from strings--
  rd<=LO;
   y<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LDY_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LDY_ZERO_PAGE_STATE_1;

when LDY_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LDY_ZERO_PAGE_STATE_2;

when LDY_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=LDY_ZERO_PAGE_STATE_3;

when LDY_ZERO_PAGE_STATE_3=> --- OPERATION

-- start from strings--
  rd<=LO;
   y<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when LDY_ZERO_PAGE_X_STATE_0=> --- OPERATION

-- start from strings--
  rd<=LO;
   y<=data;

-- end  start from strings--
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LSR_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LSR_ABSOLUTE_STATE_1;

when LSR_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LSR_ABSOLUTE_STATE_2;

when LSR_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=LSR_ABSOLUTE_STATE_3;

when LSR_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=LSR_ABSOLUTE_STATE_4;

when LSR_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=LSR_ABSOLUTE_STATE_5;

when LSR_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when LSR_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- accumulator NOT IMPLEMENTED ----
when LSR_ACCUMULATOR_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when LSR_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=LSR_ZERO_PAGE_STATE_1;

when LSR_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=LSR_ZERO_PAGE_STATE_2;

when LSR_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=LSR_ZERO_PAGE_STATE_3;

when LSR_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when LSR_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when NOP_IMPLIED_STATE_0=> --- OPERATION

-- start from strings--
    --- do nothing

-- end  start from strings--
    next_state<=NEW_INSTRUCTION;



when ORA_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ORA_ABSOLUTE_STATE_1;

when ORA_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ORA_ABSOLUTE_STATE_2;

when ORA_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=ORA_ABSOLUTE_STATE_3;

when ORA_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=ORA_ABSOLUTE_STATE_4;

when ORA_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=ORA_ABSOLUTE_STATE_5;

when ORA_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when ORA_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when ORA_ABSOLUTE_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ORA_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=ORA_IMMEDIATE_STATE_1;
when ORA_IMMEDIATE_STATE_1=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when ORA_INDIRECT_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when ORA_INDIRECT_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ORA_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ORA_ZERO_PAGE_STATE_1;

when ORA_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ORA_ZERO_PAGE_STATE_2;

when ORA_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=ORA_ZERO_PAGE_STATE_3;

when ORA_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when ORA_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when PHA_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when PHP_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when PLA_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when PLP_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- internal NOT IMPLEMENTED ----
when RESET_INTERNAL_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ROL_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ROL_ABSOLUTE_STATE_1;

when ROL_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ROL_ABSOLUTE_STATE_2;

when ROL_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=ROL_ABSOLUTE_STATE_3;

when ROL_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=ROL_ABSOLUTE_STATE_4;

when ROL_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=ROL_ABSOLUTE_STATE_5;

when ROL_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when ROL_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- accumulator NOT IMPLEMENTED ----
when ROL_ACCUMULATOR_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ROL_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ROL_ZERO_PAGE_STATE_1;

when ROL_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ROL_ZERO_PAGE_STATE_2;

when ROL_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=ROL_ZERO_PAGE_STATE_3;

when ROL_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when ROL_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ROR_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ROR_ABSOLUTE_STATE_1;

when ROR_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ROR_ABSOLUTE_STATE_2;

when ROR_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=ROR_ABSOLUTE_STATE_3;

when ROR_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=ROR_ABSOLUTE_STATE_4;

when ROR_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=ROR_ABSOLUTE_STATE_5;

when ROR_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when ROR_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- accumulator NOT IMPLEMENTED ----
when ROR_ACCUMULATOR_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when ROR_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=ROR_ZERO_PAGE_STATE_1;

when ROR_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=ROR_ZERO_PAGE_STATE_2;

when ROR_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=ROR_ZERO_PAGE_STATE_3;

when ROR_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when ROR_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when RTI_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when RTS_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;



when SBC_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=SBC_ABSOLUTE_STATE_1;

when SBC_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=SBC_ABSOLUTE_STATE_2;

when SBC_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=SBC_ABSOLUTE_STATE_3;

when SBC_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=SBC_ABSOLUTE_STATE_4;

when SBC_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=SBC_ABSOLUTE_STATE_5;

when SBC_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when SBC_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when SBC_ABSOLUTE_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when SBC_IMMEDIATE_STATE_0=>
       mem_addr<=pc_r;
       pc<=pc_r+1;
       next_state<=SBC_IMMEDIATE_STATE_1;
when SBC_IMMEDIATE_STATE_1=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when SBC_INDIRECT_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when SBC_INDIRECT_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when SBC_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=SBC_ZERO_PAGE_STATE_1;

when SBC_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=SBC_ZERO_PAGE_STATE_2;

when SBC_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=SBC_ZERO_PAGE_STATE_3;

when SBC_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when SBC_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when SEC_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when SED_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when SEI_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when STA_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=STA_ABSOLUTE_STATE_1;

when STA_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=STA_ABSOLUTE_STATE_2;

when STA_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=STA_ABSOLUTE_STATE_3;

when STA_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=STA_ABSOLUTE_STATE_4;

when STA_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=STA_ABSOLUTE_STATE_5;

when STA_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


--- absolute_y NOT IMPLEMENTED ----
when STA_ABSOLUTE_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


--- indirect_x NOT IMPLEMENTED ----
when STA_INDIRECT_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


--- indirect_y NOT IMPLEMENTED ----
when STA_INDIRECT_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;



when STA_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=STA_ZERO_PAGE_STATE_1;

when STA_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=STA_ZERO_PAGE_STATE_2;

when STA_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=STA_ZERO_PAGE_STATE_3;

when STA_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when STA_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


--- absolute_x NOT IMPLEMENTED ----
when STA_ABSOLUTE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


--- internal NOT IMPLEMENTED ----
when S_IRQ_INTERNAL_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


--- internal NOT IMPLEMENTED ----
when S_NMI_INTERNAL_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;



when STX_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=STX_ABSOLUTE_STATE_1;

when STX_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=STX_ABSOLUTE_STATE_2;

when STX_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=STX_ABSOLUTE_STATE_3;

when STX_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=STX_ABSOLUTE_STATE_4;

when STX_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=STX_ABSOLUTE_STATE_5;

when STX_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;



when STX_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=STX_ZERO_PAGE_STATE_1;

when STX_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=STX_ZERO_PAGE_STATE_2;

when STX_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=STX_ZERO_PAGE_STATE_3;

when STX_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


--- zeropage_y NOT IMPLEMENTED ----
when STX_ZERO_PAGE_Y_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;



when STY_ABSOLUTE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=STY_ABSOLUTE_STATE_1;

when STY_ABSOLUTE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=STY_ABSOLUTE_STATE_2;

when STY_ABSOLUTE_STATE_2=>
     mem_addr<=mem_addr_r+1;
     next_state<=STY_ABSOLUTE_STATE_3;

when STY_ABSOLUTE_STATE_3=>
    rd<=LO;
      addr_hi<=data;
      next_state<=STY_ABSOLUTE_STATE_4;

when STY_ABSOLUTE_STATE_4=>
     mem_addr<=addr_hi_r&addr_lo_r;
     pc<=pc_r+2;
     next_state<=STY_ABSOLUTE_STATE_5;

when STY_ABSOLUTE_STATE_5=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;



when STY_ZERO_PAGE_STATE_0=>
       mem_addr<=pc_r;
       next_state<=STY_ZERO_PAGE_STATE_1;

when STY_ZERO_PAGE_STATE_1=>
    rd<=LO;
    addr_lo<=data;
    next_state<=STY_ZERO_PAGE_STATE_2;

when STY_ZERO_PAGE_STATE_2=>
     mem_addr<="00000000" & addr_lo_r;
     pc<=pc_r+1;
     next_state<=STY_ZERO_PAGE_STATE_3;

when STY_ZERO_PAGE_STATE_3=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---zeropagex NOT IMPLEMENTED ----
when STY_ZERO_PAGE_X_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when TAX_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when TAY_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when TSX_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when TXA_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
--- NOT IMPLEMENTED ----
--- NOT IMPLEMENTED ----
    next_state<=NEW_INSTRUCTION;


---  implied NOT IMPLEMENTED ----
when TXS_IMPLIED_STATE_0=> --- OPERATION
----- NOT IMPLEMENTED (no string)
    next_state<=NEW_INSTRUCTION;
when others=>
next_state<=NEW_INSTRUCTION;
end case;
end process;
end c6502_architecture;
